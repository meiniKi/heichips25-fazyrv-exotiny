module heichips25_fazyrv_exotiny (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire ccx_req;
 wire gpo;
 wire \i_exotiny._0000_ ;
 wire \i_exotiny._0013_[0] ;
 wire \i_exotiny._0013_[1] ;
 wire \i_exotiny._0013_[2] ;
 wire \i_exotiny._0013_[3] ;
 wire \i_exotiny._0014_[0] ;
 wire \i_exotiny._0014_[1] ;
 wire \i_exotiny._0014_[2] ;
 wire \i_exotiny._0014_[3] ;
 wire \i_exotiny._0015_[0] ;
 wire \i_exotiny._0015_[1] ;
 wire \i_exotiny._0015_[2] ;
 wire \i_exotiny._0015_[3] ;
 wire \i_exotiny._0016_[0] ;
 wire \i_exotiny._0016_[1] ;
 wire \i_exotiny._0016_[2] ;
 wire \i_exotiny._0016_[3] ;
 wire \i_exotiny._0017_[0] ;
 wire \i_exotiny._0017_[1] ;
 wire \i_exotiny._0017_[2] ;
 wire \i_exotiny._0017_[3] ;
 wire \i_exotiny._0018_[0] ;
 wire \i_exotiny._0018_[1] ;
 wire \i_exotiny._0018_[2] ;
 wire \i_exotiny._0018_[3] ;
 wire \i_exotiny._0019_[0] ;
 wire \i_exotiny._0019_[1] ;
 wire \i_exotiny._0019_[2] ;
 wire \i_exotiny._0019_[3] ;
 wire \i_exotiny._0020_[0] ;
 wire \i_exotiny._0020_[1] ;
 wire \i_exotiny._0020_[2] ;
 wire \i_exotiny._0020_[3] ;
 wire \i_exotiny._0021_[0] ;
 wire \i_exotiny._0021_[1] ;
 wire \i_exotiny._0021_[2] ;
 wire \i_exotiny._0021_[3] ;
 wire \i_exotiny._0022_[0] ;
 wire \i_exotiny._0022_[1] ;
 wire \i_exotiny._0022_[2] ;
 wire \i_exotiny._0022_[3] ;
 wire \i_exotiny._0023_[0] ;
 wire \i_exotiny._0023_[1] ;
 wire \i_exotiny._0023_[2] ;
 wire \i_exotiny._0023_[3] ;
 wire \i_exotiny._0024_[0] ;
 wire \i_exotiny._0024_[1] ;
 wire \i_exotiny._0024_[2] ;
 wire \i_exotiny._0024_[3] ;
 wire \i_exotiny._0025_[0] ;
 wire \i_exotiny._0025_[1] ;
 wire \i_exotiny._0025_[2] ;
 wire \i_exotiny._0025_[3] ;
 wire \i_exotiny._0026_[0] ;
 wire \i_exotiny._0026_[1] ;
 wire \i_exotiny._0026_[2] ;
 wire \i_exotiny._0026_[3] ;
 wire \i_exotiny._0027_[0] ;
 wire \i_exotiny._0027_[1] ;
 wire \i_exotiny._0027_[2] ;
 wire \i_exotiny._0027_[3] ;
 wire \i_exotiny._0028_[0] ;
 wire \i_exotiny._0028_[1] ;
 wire \i_exotiny._0028_[2] ;
 wire \i_exotiny._0028_[3] ;
 wire \i_exotiny._0029_[0] ;
 wire \i_exotiny._0029_[1] ;
 wire \i_exotiny._0029_[2] ;
 wire \i_exotiny._0029_[3] ;
 wire \i_exotiny._0030_[0] ;
 wire \i_exotiny._0030_[1] ;
 wire \i_exotiny._0030_[2] ;
 wire \i_exotiny._0030_[3] ;
 wire \i_exotiny._0031_[0] ;
 wire \i_exotiny._0031_[1] ;
 wire \i_exotiny._0031_[2] ;
 wire \i_exotiny._0031_[3] ;
 wire \i_exotiny._0032_[0] ;
 wire \i_exotiny._0032_[1] ;
 wire \i_exotiny._0032_[2] ;
 wire \i_exotiny._0032_[3] ;
 wire \i_exotiny._0033_[0] ;
 wire \i_exotiny._0033_[1] ;
 wire \i_exotiny._0033_[2] ;
 wire \i_exotiny._0033_[3] ;
 wire \i_exotiny._0034_[0] ;
 wire \i_exotiny._0034_[1] ;
 wire \i_exotiny._0034_[2] ;
 wire \i_exotiny._0034_[3] ;
 wire \i_exotiny._0035_[0] ;
 wire \i_exotiny._0035_[1] ;
 wire \i_exotiny._0035_[2] ;
 wire \i_exotiny._0035_[3] ;
 wire \i_exotiny._0036_[0] ;
 wire \i_exotiny._0036_[1] ;
 wire \i_exotiny._0036_[2] ;
 wire \i_exotiny._0036_[3] ;
 wire \i_exotiny._0037_[0] ;
 wire \i_exotiny._0037_[1] ;
 wire \i_exotiny._0037_[2] ;
 wire \i_exotiny._0037_[3] ;
 wire \i_exotiny._0038_[0] ;
 wire \i_exotiny._0038_[1] ;
 wire \i_exotiny._0038_[2] ;
 wire \i_exotiny._0038_[3] ;
 wire \i_exotiny._0039_[0] ;
 wire \i_exotiny._0039_[1] ;
 wire \i_exotiny._0039_[2] ;
 wire \i_exotiny._0039_[3] ;
 wire \i_exotiny._0040_[0] ;
 wire \i_exotiny._0040_[1] ;
 wire \i_exotiny._0040_[2] ;
 wire \i_exotiny._0040_[3] ;
 wire \i_exotiny._0041_[0] ;
 wire \i_exotiny._0041_[1] ;
 wire \i_exotiny._0041_[2] ;
 wire \i_exotiny._0041_[3] ;
 wire \i_exotiny._0042_[0] ;
 wire \i_exotiny._0042_[1] ;
 wire \i_exotiny._0042_[2] ;
 wire \i_exotiny._0042_[3] ;
 wire \i_exotiny._0043_[0] ;
 wire \i_exotiny._0043_[1] ;
 wire \i_exotiny._0043_[2] ;
 wire \i_exotiny._0043_[3] ;
 wire \i_exotiny._0077_[0] ;
 wire \i_exotiny._0077_[1] ;
 wire \i_exotiny._0077_[2] ;
 wire \i_exotiny._0077_[3] ;
 wire \i_exotiny._0077_[4] ;
 wire \i_exotiny._0079_[0] ;
 wire \i_exotiny._0079_[1] ;
 wire \i_exotiny._0079_[2] ;
 wire \i_exotiny._0079_[3] ;
 wire \i_exotiny._0079_[4] ;
 wire \i_exotiny._0314_[10] ;
 wire \i_exotiny._0314_[11] ;
 wire \i_exotiny._0314_[12] ;
 wire \i_exotiny._0314_[13] ;
 wire \i_exotiny._0314_[14] ;
 wire \i_exotiny._0314_[15] ;
 wire \i_exotiny._0314_[16] ;
 wire \i_exotiny._0314_[17] ;
 wire \i_exotiny._0314_[18] ;
 wire \i_exotiny._0314_[19] ;
 wire \i_exotiny._0314_[20] ;
 wire \i_exotiny._0314_[21] ;
 wire \i_exotiny._0314_[22] ;
 wire \i_exotiny._0314_[23] ;
 wire \i_exotiny._0314_[24] ;
 wire \i_exotiny._0314_[25] ;
 wire \i_exotiny._0314_[26] ;
 wire \i_exotiny._0314_[27] ;
 wire \i_exotiny._0314_[28] ;
 wire \i_exotiny._0314_[29] ;
 wire \i_exotiny._0314_[2] ;
 wire \i_exotiny._0314_[30] ;
 wire \i_exotiny._0314_[31] ;
 wire \i_exotiny._0314_[3] ;
 wire \i_exotiny._0314_[4] ;
 wire \i_exotiny._0314_[5] ;
 wire \i_exotiny._0314_[6] ;
 wire \i_exotiny._0314_[7] ;
 wire \i_exotiny._0314_[8] ;
 wire \i_exotiny._0314_[9] ;
 wire \i_exotiny._0315_[10] ;
 wire \i_exotiny._0315_[11] ;
 wire \i_exotiny._0315_[12] ;
 wire \i_exotiny._0315_[13] ;
 wire \i_exotiny._0315_[14] ;
 wire \i_exotiny._0315_[15] ;
 wire \i_exotiny._0315_[16] ;
 wire \i_exotiny._0315_[17] ;
 wire \i_exotiny._0315_[18] ;
 wire \i_exotiny._0315_[19] ;
 wire \i_exotiny._0315_[20] ;
 wire \i_exotiny._0315_[21] ;
 wire \i_exotiny._0315_[22] ;
 wire \i_exotiny._0315_[23] ;
 wire \i_exotiny._0315_[24] ;
 wire \i_exotiny._0315_[25] ;
 wire \i_exotiny._0315_[26] ;
 wire \i_exotiny._0315_[27] ;
 wire \i_exotiny._0315_[28] ;
 wire \i_exotiny._0315_[29] ;
 wire \i_exotiny._0315_[2] ;
 wire \i_exotiny._0315_[30] ;
 wire \i_exotiny._0315_[31] ;
 wire \i_exotiny._0315_[3] ;
 wire \i_exotiny._0315_[4] ;
 wire \i_exotiny._0315_[5] ;
 wire \i_exotiny._0315_[6] ;
 wire \i_exotiny._0315_[7] ;
 wire \i_exotiny._0315_[8] ;
 wire \i_exotiny._0315_[9] ;
 wire \i_exotiny._0327_[0] ;
 wire \i_exotiny._0327_[1] ;
 wire \i_exotiny._0352_ ;
 wire \i_exotiny._0369_[0] ;
 wire \i_exotiny._0369_[10] ;
 wire \i_exotiny._0369_[11] ;
 wire \i_exotiny._0369_[12] ;
 wire \i_exotiny._0369_[13] ;
 wire \i_exotiny._0369_[14] ;
 wire \i_exotiny._0369_[15] ;
 wire \i_exotiny._0369_[16] ;
 wire \i_exotiny._0369_[17] ;
 wire \i_exotiny._0369_[18] ;
 wire \i_exotiny._0369_[19] ;
 wire \i_exotiny._0369_[1] ;
 wire \i_exotiny._0369_[20] ;
 wire \i_exotiny._0369_[21] ;
 wire \i_exotiny._0369_[22] ;
 wire \i_exotiny._0369_[23] ;
 wire \i_exotiny._0369_[24] ;
 wire \i_exotiny._0369_[25] ;
 wire \i_exotiny._0369_[26] ;
 wire \i_exotiny._0369_[27] ;
 wire \i_exotiny._0369_[28] ;
 wire \i_exotiny._0369_[29] ;
 wire \i_exotiny._0369_[2] ;
 wire \i_exotiny._0369_[30] ;
 wire \i_exotiny._0369_[3] ;
 wire \i_exotiny._0369_[4] ;
 wire \i_exotiny._0369_[5] ;
 wire \i_exotiny._0369_[6] ;
 wire \i_exotiny._0369_[7] ;
 wire \i_exotiny._0369_[8] ;
 wire \i_exotiny._0369_[9] ;
 wire \i_exotiny._0542_ ;
 wire \i_exotiny._0550_ ;
 wire \i_exotiny._0571_ ;
 wire \i_exotiny._0590_ ;
 wire \i_exotiny._0601_ ;
 wire \i_exotiny._1160_[0] ;
 wire \i_exotiny._1160_[10] ;
 wire \i_exotiny._1160_[11] ;
 wire \i_exotiny._1160_[12] ;
 wire \i_exotiny._1160_[13] ;
 wire \i_exotiny._1160_[14] ;
 wire \i_exotiny._1160_[15] ;
 wire \i_exotiny._1160_[16] ;
 wire \i_exotiny._1160_[17] ;
 wire \i_exotiny._1160_[18] ;
 wire \i_exotiny._1160_[19] ;
 wire \i_exotiny._1160_[1] ;
 wire \i_exotiny._1160_[20] ;
 wire \i_exotiny._1160_[21] ;
 wire \i_exotiny._1160_[22] ;
 wire \i_exotiny._1160_[23] ;
 wire \i_exotiny._1160_[24] ;
 wire \i_exotiny._1160_[25] ;
 wire \i_exotiny._1160_[26] ;
 wire \i_exotiny._1160_[27] ;
 wire \i_exotiny._1160_[2] ;
 wire \i_exotiny._1160_[3] ;
 wire \i_exotiny._1160_[4] ;
 wire \i_exotiny._1160_[5] ;
 wire \i_exotiny._1160_[6] ;
 wire \i_exotiny._1160_[7] ;
 wire \i_exotiny._1160_[8] ;
 wire \i_exotiny._1160_[9] ;
 wire \i_exotiny._1206_ ;
 wire \i_exotiny._1207_ ;
 wire \i_exotiny._1265_ ;
 wire \i_exotiny._1266_ ;
 wire \i_exotiny._1306_ ;
 wire \i_exotiny._1308_ ;
 wire \i_exotiny._1309_ ;
 wire \i_exotiny._1311_ ;
 wire \i_exotiny._1312_ ;
 wire \i_exotiny._1429_ ;
 wire \i_exotiny._1465_ ;
 wire \i_exotiny._1489_[0] ;
 wire \i_exotiny._1489_[1] ;
 wire \i_exotiny._1489_[2] ;
 wire \i_exotiny._1489_[3] ;
 wire \i_exotiny._1586_ ;
 wire \i_exotiny._1611_[10] ;
 wire \i_exotiny._1611_[11] ;
 wire \i_exotiny._1611_[13] ;
 wire \i_exotiny._1611_[14] ;
 wire \i_exotiny._1611_[15] ;
 wire \i_exotiny._1611_[17] ;
 wire \i_exotiny._1611_[18] ;
 wire \i_exotiny._1611_[19] ;
 wire \i_exotiny._1611_[1] ;
 wire \i_exotiny._1611_[21] ;
 wire \i_exotiny._1611_[22] ;
 wire \i_exotiny._1611_[23] ;
 wire \i_exotiny._1611_[25] ;
 wire \i_exotiny._1611_[26] ;
 wire \i_exotiny._1611_[27] ;
 wire \i_exotiny._1611_[29] ;
 wire \i_exotiny._1611_[2] ;
 wire \i_exotiny._1611_[30] ;
 wire \i_exotiny._1611_[31] ;
 wire \i_exotiny._1611_[3] ;
 wire \i_exotiny._1611_[5] ;
 wire \i_exotiny._1611_[6] ;
 wire \i_exotiny._1611_[7] ;
 wire \i_exotiny._1611_[9] ;
 wire \i_exotiny._1612_[0] ;
 wire \i_exotiny._1612_[1] ;
 wire \i_exotiny._1612_[2] ;
 wire \i_exotiny._1612_[3] ;
 wire \i_exotiny._1614_[0] ;
 wire \i_exotiny._1614_[1] ;
 wire \i_exotiny._1614_[2] ;
 wire \i_exotiny._1614_[3] ;
 wire \i_exotiny._1615_[0] ;
 wire \i_exotiny._1615_[1] ;
 wire \i_exotiny._1615_[2] ;
 wire \i_exotiny._1615_[3] ;
 wire \i_exotiny._1616_[0] ;
 wire \i_exotiny._1616_[1] ;
 wire \i_exotiny._1616_[2] ;
 wire \i_exotiny._1616_[3] ;
 wire \i_exotiny._1617_[0] ;
 wire \i_exotiny._1617_[1] ;
 wire \i_exotiny._1617_[2] ;
 wire \i_exotiny._1617_[3] ;
 wire \i_exotiny._1618_[0] ;
 wire \i_exotiny._1618_[1] ;
 wire \i_exotiny._1618_[2] ;
 wire \i_exotiny._1618_[3] ;
 wire \i_exotiny._1619_[0] ;
 wire \i_exotiny._1619_[1] ;
 wire \i_exotiny._1619_[2] ;
 wire \i_exotiny._1619_[3] ;
 wire \i_exotiny._1623_ ;
 wire \i_exotiny._1652_[0] ;
 wire \i_exotiny._1660_ ;
 wire clk_regs;
 wire \i_exotiny._1711_ ;
 wire \i_exotiny._1715_ ;
 wire \i_exotiny._1725_ ;
 wire \i_exotiny._1737_ ;
 wire \i_exotiny._1757_ ;
 wire \i_exotiny._1793_ ;
 wire \i_exotiny._1840_[11] ;
 wire \i_exotiny._1902_[0] ;
 wire \i_exotiny._1902_[1] ;
 wire \i_exotiny._1902_[2] ;
 wire \i_exotiny._1902_[3] ;
 wire \i_exotiny._1902_[4] ;
 wire \i_exotiny._1902_[5] ;
 wire \i_exotiny._1902_[6] ;
 wire \i_exotiny._1924_[10] ;
 wire \i_exotiny._1924_[11] ;
 wire \i_exotiny._1924_[12] ;
 wire \i_exotiny._1924_[13] ;
 wire \i_exotiny._1924_[14] ;
 wire \i_exotiny._1924_[15] ;
 wire \i_exotiny._1924_[16] ;
 wire \i_exotiny._1924_[17] ;
 wire \i_exotiny._1924_[18] ;
 wire \i_exotiny._1924_[19] ;
 wire \i_exotiny._1924_[1] ;
 wire \i_exotiny._1924_[20] ;
 wire \i_exotiny._1924_[21] ;
 wire \i_exotiny._1924_[22] ;
 wire \i_exotiny._1924_[23] ;
 wire \i_exotiny._1924_[24] ;
 wire \i_exotiny._1924_[25] ;
 wire \i_exotiny._1924_[26] ;
 wire \i_exotiny._1924_[27] ;
 wire \i_exotiny._1924_[28] ;
 wire \i_exotiny._1924_[29] ;
 wire \i_exotiny._1924_[2] ;
 wire \i_exotiny._1924_[30] ;
 wire \i_exotiny._1924_[31] ;
 wire \i_exotiny._1924_[3] ;
 wire \i_exotiny._1924_[4] ;
 wire \i_exotiny._1924_[5] ;
 wire \i_exotiny._1924_[6] ;
 wire \i_exotiny._1924_[7] ;
 wire \i_exotiny._1924_[8] ;
 wire \i_exotiny._1924_[9] ;
 wire \i_exotiny._1956_ ;
 wire \i_exotiny._2025_[3] ;
 wire \i_exotiny._2025_[4] ;
 wire \i_exotiny._2025_[5] ;
 wire \i_exotiny._2025_[6] ;
 wire \i_exotiny._2032_ ;
 wire \i_exotiny._2034_[0] ;
 wire \i_exotiny._2034_[1] ;
 wire \i_exotiny._2034_[2] ;
 wire \i_exotiny._2034_[3] ;
 wire \i_exotiny._2034_[4] ;
 wire \i_exotiny._2034_[5] ;
 wire \i_exotiny._2034_[6] ;
 wire \i_exotiny._2034_[7] ;
 wire \i_exotiny._2034_[8] ;
 wire \i_exotiny._2034_[9] ;
 wire \i_exotiny._2043_[0] ;
 wire \i_exotiny._2043_[1] ;
 wire \i_exotiny._2043_[2] ;
 wire \i_exotiny._2043_[3] ;
 wire \i_exotiny._2043_[4] ;
 wire \i_exotiny._2043_[5] ;
 wire \i_exotiny._2043_[6] ;
 wire \i_exotiny._2043_[7] ;
 wire \i_exotiny._2043_[8] ;
 wire \i_exotiny._2043_[9] ;
 wire \i_exotiny._2044_[1] ;
 wire \i_exotiny._2055_[0] ;
 wire \i_exotiny._2055_[1] ;
 wire \i_exotiny._2055_[2] ;
 wire \i_exotiny._2160_ ;
 wire \i_exotiny._3871_ ;
 wire \i_exotiny._6090_[0] ;
 wire \i_exotiny._6090_[1] ;
 wire \i_exotiny._6090_[2] ;
 wire \i_exotiny._6090_[3] ;
 wire \i_exotiny.core_res_en_n ;
 wire \i_exotiny.gpo[0] ;
 wire \i_exotiny.gpo[1] ;
 wire \i_exotiny.gpo[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[10] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[11] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[12] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[13] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[14] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[15] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[16] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[17] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[18] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[19] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[20] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[21] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[22] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[23] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[24] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[25] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[26] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[27] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[28] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[29] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[30] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[31] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[4] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[5] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[6] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[7] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[8] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[9] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ;
 wire \i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_hlt_pc_ccx ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[4] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[5] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[2] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[3] ;
 wire \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r ;
 wire \i_exotiny.i_rstctl.cnt[0] ;
 wire \i_exotiny.i_rstctl.cnt[1] ;
 wire \i_exotiny.i_rstctl.cnt[2] ;
 wire \i_exotiny.i_rstctl.cnt[3] ;
 wire \i_exotiny.i_rstctl.cnt[4] ;
 wire \i_exotiny.i_rstctl.cnt[5] ;
 wire \i_exotiny.i_rstctl.cnt[6] ;
 wire \i_exotiny.i_rstctl.sys_res_n ;
 wire \i_exotiny.i_rstctl.wdg_res_n ;
 wire \i_exotiny.i_wb_qspi_mem.cnt_r[1] ;
 wire \i_exotiny.i_wb_qspi_mem.cnt_r[2] ;
 wire \i_exotiny.i_wb_qspi_mem.crm_r ;
 wire \i_exotiny.i_wb_regs.spi_auto_cs_o ;
 wire \i_exotiny.i_wb_regs.spi_cpol_o ;
 wire \i_exotiny.i_wb_regs.spi_size_o[0] ;
 wire \i_exotiny.i_wb_regs.spi_size_o[1] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[1] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[2] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[3] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[4] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[5] ;
 wire \i_exotiny.i_wb_spi.cnt_hbit_r[6] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[0] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[1] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[2] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[3] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[4] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[5] ;
 wire \i_exotiny.i_wb_spi.cnt_presc_r[6] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[0] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[10] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[11] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[12] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[13] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[14] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[15] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[16] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[17] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[18] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[19] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[1] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[20] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[21] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[22] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[23] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[24] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[25] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[26] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[27] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[28] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[29] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[2] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[30] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[31] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[3] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[4] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[5] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[6] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[7] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[8] ;
 wire \i_exotiny.i_wb_spi.dat_rx_r[9] ;
 wire \i_exotiny.i_wb_spi.sck_r ;
 wire \i_exotiny.i_wb_spi.spi_sdo_o ;
 wire \i_exotiny.i_wb_spi.state_r[0] ;
 wire \i_exotiny.i_wb_spi.state_r[10] ;
 wire \i_exotiny.i_wb_spi.state_r[11] ;
 wire \i_exotiny.i_wb_spi.state_r[12] ;
 wire \i_exotiny.i_wb_spi.state_r[13] ;
 wire \i_exotiny.i_wb_spi.state_r[14] ;
 wire \i_exotiny.i_wb_spi.state_r[15] ;
 wire \i_exotiny.i_wb_spi.state_r[16] ;
 wire \i_exotiny.i_wb_spi.state_r[17] ;
 wire \i_exotiny.i_wb_spi.state_r[18] ;
 wire \i_exotiny.i_wb_spi.state_r[19] ;
 wire \i_exotiny.i_wb_spi.state_r[1] ;
 wire \i_exotiny.i_wb_spi.state_r[20] ;
 wire \i_exotiny.i_wb_spi.state_r[21] ;
 wire \i_exotiny.i_wb_spi.state_r[22] ;
 wire \i_exotiny.i_wb_spi.state_r[23] ;
 wire \i_exotiny.i_wb_spi.state_r[24] ;
 wire \i_exotiny.i_wb_spi.state_r[25] ;
 wire \i_exotiny.i_wb_spi.state_r[26] ;
 wire \i_exotiny.i_wb_spi.state_r[27] ;
 wire \i_exotiny.i_wb_spi.state_r[28] ;
 wire \i_exotiny.i_wb_spi.state_r[29] ;
 wire \i_exotiny.i_wb_spi.state_r[2] ;
 wire \i_exotiny.i_wb_spi.state_r[30] ;
 wire \i_exotiny.i_wb_spi.state_r[31] ;
 wire \i_exotiny.i_wb_spi.state_r[3] ;
 wire \i_exotiny.i_wb_spi.state_r[4] ;
 wire \i_exotiny.i_wb_spi.state_r[5] ;
 wire \i_exotiny.i_wb_spi.state_r[6] ;
 wire \i_exotiny.i_wb_spi.state_r[7] ;
 wire \i_exotiny.i_wb_spi.state_r[8] ;
 wire \i_exotiny.i_wb_spi.state_r[9] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[0] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[10] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[11] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[12] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[13] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[14] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[15] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[16] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[17] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[18] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[19] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[1] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[2] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[3] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[4] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[5] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[6] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[7] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[8] ;
 wire \i_exotiny.i_wdg_top.clk_div_inst.cnt[9] ;
 wire \i_exotiny.i_wdg_top.cntr_inst.rst_n_sync ;
 wire \i_exotiny.i_wdg_top.do_cnt ;
 wire \i_exotiny.i_wdg_top.fsm_inst.sw_trg_s1wto ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[0] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[10] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[11] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[12] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[13] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[1] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[2] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[3] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[4] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[5] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[6] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[7] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[8] ;
 wire \i_exotiny.i_wdg_top.o_wb_dat[9] ;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net42;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_57_clk_regs;
 wire clknet_leaf_58_clk_regs;
 wire clknet_leaf_59_clk_regs;
 wire clknet_leaf_60_clk_regs;
 wire clknet_leaf_61_clk_regs;
 wire clknet_leaf_62_clk_regs;
 wire clknet_leaf_63_clk_regs;
 wire clknet_leaf_64_clk_regs;
 wire clknet_leaf_65_clk_regs;
 wire clknet_leaf_66_clk_regs;
 wire clknet_leaf_67_clk_regs;
 wire clknet_leaf_68_clk_regs;
 wire clknet_leaf_69_clk_regs;
 wire clknet_leaf_70_clk_regs;
 wire clknet_leaf_71_clk_regs;
 wire clknet_leaf_72_clk_regs;
 wire clknet_leaf_73_clk_regs;
 wire clknet_leaf_74_clk_regs;
 wire clknet_leaf_75_clk_regs;
 wire clknet_leaf_76_clk_regs;
 wire clknet_leaf_77_clk_regs;
 wire clknet_leaf_78_clk_regs;
 wire clknet_leaf_79_clk_regs;
 wire clknet_leaf_80_clk_regs;
 wire clknet_leaf_81_clk_regs;
 wire clknet_leaf_82_clk_regs;
 wire clknet_leaf_83_clk_regs;
 wire clknet_leaf_84_clk_regs;
 wire clknet_leaf_85_clk_regs;
 wire clknet_leaf_86_clk_regs;
 wire clknet_leaf_87_clk_regs;
 wire clknet_leaf_89_clk_regs;
 wire clknet_leaf_90_clk_regs;
 wire clknet_leaf_91_clk_regs;
 wire clknet_leaf_92_clk_regs;
 wire clknet_leaf_93_clk_regs;
 wire clknet_leaf_94_clk_regs;
 wire clknet_leaf_95_clk_regs;
 wire clknet_leaf_96_clk_regs;
 wire clknet_leaf_97_clk_regs;
 wire clknet_leaf_98_clk_regs;
 wire clknet_leaf_99_clk_regs;
 wire clknet_leaf_100_clk_regs;
 wire clknet_leaf_101_clk_regs;
 wire clknet_leaf_102_clk_regs;
 wire clknet_leaf_103_clk_regs;
 wire clknet_leaf_104_clk_regs;
 wire clknet_leaf_105_clk_regs;
 wire clknet_leaf_106_clk_regs;
 wire clknet_leaf_107_clk_regs;
 wire clknet_leaf_108_clk_regs;
 wire clknet_leaf_109_clk_regs;
 wire clknet_leaf_110_clk_regs;
 wire clknet_leaf_111_clk_regs;
 wire clknet_leaf_112_clk_regs;
 wire clknet_leaf_113_clk_regs;
 wire clknet_leaf_114_clk_regs;
 wire clknet_leaf_115_clk_regs;
 wire clknet_leaf_116_clk_regs;
 wire clknet_leaf_117_clk_regs;
 wire clknet_leaf_118_clk_regs;
 wire clknet_leaf_119_clk_regs;
 wire clknet_leaf_120_clk_regs;
 wire clknet_leaf_121_clk_regs;
 wire clknet_leaf_122_clk_regs;
 wire clknet_leaf_123_clk_regs;
 wire clknet_leaf_124_clk_regs;
 wire clknet_leaf_125_clk_regs;
 wire clknet_leaf_126_clk_regs;
 wire clknet_leaf_127_clk_regs;
 wire clknet_leaf_128_clk_regs;
 wire clknet_leaf_129_clk_regs;
 wire clknet_leaf_130_clk_regs;
 wire clknet_leaf_131_clk_regs;
 wire clknet_leaf_132_clk_regs;
 wire clknet_leaf_133_clk_regs;
 wire clknet_leaf_134_clk_regs;
 wire clknet_leaf_135_clk_regs;
 wire clknet_leaf_136_clk_regs;
 wire clknet_leaf_137_clk_regs;
 wire clknet_leaf_138_clk_regs;
 wire clknet_leaf_139_clk_regs;
 wire clknet_leaf_140_clk_regs;
 wire clknet_leaf_141_clk_regs;
 wire clknet_leaf_142_clk_regs;
 wire clknet_leaf_143_clk_regs;
 wire clknet_leaf_144_clk_regs;
 wire clknet_leaf_145_clk_regs;
 wire clknet_leaf_146_clk_regs;
 wire clknet_leaf_147_clk_regs;
 wire clknet_leaf_148_clk_regs;
 wire clknet_leaf_149_clk_regs;
 wire clknet_leaf_150_clk_regs;
 wire clknet_leaf_151_clk_regs;
 wire clknet_leaf_152_clk_regs;
 wire clknet_leaf_153_clk_regs;
 wire clknet_leaf_154_clk_regs;
 wire clknet_leaf_155_clk_regs;
 wire clknet_leaf_156_clk_regs;
 wire clknet_leaf_157_clk_regs;
 wire clknet_leaf_158_clk_regs;
 wire clknet_leaf_159_clk_regs;
 wire clknet_leaf_160_clk_regs;
 wire clknet_leaf_161_clk_regs;
 wire clknet_leaf_162_clk_regs;
 wire clknet_leaf_163_clk_regs;
 wire clknet_leaf_164_clk_regs;
 wire clknet_leaf_165_clk_regs;
 wire clknet_leaf_166_clk_regs;
 wire clknet_leaf_167_clk_regs;
 wire clknet_leaf_168_clk_regs;
 wire clknet_leaf_169_clk_regs;
 wire clknet_leaf_170_clk_regs;
 wire clknet_leaf_171_clk_regs;
 wire clknet_leaf_172_clk_regs;
 wire clknet_leaf_173_clk_regs;
 wire clknet_leaf_174_clk_regs;
 wire clknet_leaf_175_clk_regs;
 wire clknet_leaf_176_clk_regs;
 wire clknet_leaf_177_clk_regs;
 wire clknet_leaf_178_clk_regs;
 wire clknet_leaf_179_clk_regs;
 wire clknet_leaf_180_clk_regs;
 wire clknet_leaf_181_clk_regs;
 wire clknet_leaf_182_clk_regs;
 wire clknet_leaf_183_clk_regs;
 wire clknet_leaf_184_clk_regs;
 wire clknet_leaf_185_clk_regs;
 wire clknet_leaf_186_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire [0:0] \i_exotiny._5416_$func$/home/user/heichips25-fazyrv-exotiny/build/exotiny_preproc.v:7385$12.$result ;
 wire [0:0] \i_exotiny._5420_$func$/home/user/heichips25-fazyrv-exotiny/build/exotiny_preproc.v:7404$13.$result ;
 wire [0:0] \i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r ;
 wire [0:0] \i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data ;
 wire [0:0] \i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.genblk7.g_value.r_value ;
 wire [0:0] \i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_hw_set ;
 wire [0:0] \i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data ;
 wire [0:0] \i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.genblk7.g_value.r_value ;
 wire [0:0] \i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set ;
 wire [0:0] \i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data ;
 wire [0:0] \i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.genblk7.g_value.r_value ;
 wire [0:0] \i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data ;

 sg13g2_inv_4 _04599_ (.A(net3567),
    .Y(_01361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _04600_ (.Y(_01362_),
    .A(net3834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04601_ (.VDD(VPWR),
    .Y(_01363_),
    .A(net3824),
    .VSS(VGND));
 sg13g2_inv_1 _04602_ (.VDD(VPWR),
    .Y(_01364_),
    .A(\i_exotiny.gpo[2] ),
    .VSS(VGND));
 sg13g2_inv_4 _04603_ (.A(net3730),
    .Y(_01365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _04604_ (.A(net3624),
    .Y(_01366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04605_ (.VDD(VPWR),
    .Y(_01367_),
    .A(\i_exotiny._1615_[1] ),
    .VSS(VGND));
 sg13g2_inv_1 _04606_ (.VDD(VPWR),
    .Y(_01368_),
    .A(net3466),
    .VSS(VGND));
 sg13g2_inv_1 _04607_ (.VDD(VPWR),
    .Y(_01369_),
    .A(net2037),
    .VSS(VGND));
 sg13g2_inv_2 _04608_ (.Y(_01370_),
    .A(net2886),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _04609_ (.Y(_01371_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04610_ (.VDD(VPWR),
    .Y(_01372_),
    .A(_00019_),
    .VSS(VGND));
 sg13g2_inv_1 _04611_ (.VDD(VPWR),
    .Y(_01373_),
    .A(_00018_),
    .VSS(VGND));
 sg13g2_inv_1 _04612_ (.VDD(VPWR),
    .Y(_01374_),
    .A(_00017_),
    .VSS(VGND));
 sg13g2_inv_1 _04613_ (.VDD(VPWR),
    .Y(_01375_),
    .A(_00016_),
    .VSS(VGND));
 sg13g2_inv_1 _04614_ (.VDD(VPWR),
    .Y(_01376_),
    .A(_00015_),
    .VSS(VGND));
 sg13g2_inv_1 _04615_ (.VDD(VPWR),
    .Y(_01377_),
    .A(net3511),
    .VSS(VGND));
 sg13g2_inv_1 _04616_ (.VDD(VPWR),
    .Y(_01378_),
    .A(net1291),
    .VSS(VGND));
 sg13g2_inv_1 _04617_ (.VDD(VPWR),
    .Y(_01379_),
    .A(net3634),
    .VSS(VGND));
 sg13g2_inv_1 _04618_ (.VDD(VPWR),
    .Y(_01380_),
    .A(net1270),
    .VSS(VGND));
 sg13g2_inv_1 _04619_ (.VDD(VPWR),
    .Y(_01381_),
    .A(net3726),
    .VSS(VGND));
 sg13g2_inv_1 _04620_ (.VDD(VPWR),
    .Y(_01382_),
    .A(net1244),
    .VSS(VGND));
 sg13g2_inv_2 _04621_ (.Y(_01383_),
    .A(net1230),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _04622_ (.Y(_01384_),
    .A(net1232),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _04623_ (.A(net1267),
    .Y(_01385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _04624_ (.Y(_01386_),
    .A(net3822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04625_ (.VDD(VPWR),
    .Y(_01387_),
    .A(net3789),
    .VSS(VGND));
 sg13g2_inv_4 _04626_ (.A(net1268),
    .Y(_01388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04627_ (.VDD(VPWR),
    .Y(_01389_),
    .A(net3586),
    .VSS(VGND));
 sg13g2_inv_4 _04628_ (.A(net3762),
    .Y(_01390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _04629_ (.A(net3820),
    .Y(_01391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04630_ (.VDD(VPWR),
    .Y(_01392_),
    .A(net3788),
    .VSS(VGND));
 sg13g2_inv_4 _04631_ (.A(net3784),
    .Y(_01393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _04632_ (.Y(_01394_),
    .A(net1257),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04633_ (.VDD(VPWR),
    .Y(_01395_),
    .A(net1237),
    .VSS(VGND));
 sg13g2_inv_1 _04634_ (.VDD(VPWR),
    .Y(_01396_),
    .A(net3838),
    .VSS(VGND));
 sg13g2_inv_1 _04635_ (.VDD(VPWR),
    .Y(_01397_),
    .A(net1961),
    .VSS(VGND));
 sg13g2_inv_1 _04636_ (.VDD(VPWR),
    .Y(_01398_),
    .A(\i_exotiny._2034_[0] ),
    .VSS(VGND));
 sg13g2_inv_1 _04637_ (.VDD(VPWR),
    .Y(_01399_),
    .A(\i_exotiny._2034_[1] ),
    .VSS(VGND));
 sg13g2_inv_1 _04638_ (.VDD(VPWR),
    .Y(_01400_),
    .A(\i_exotiny._2034_[2] ),
    .VSS(VGND));
 sg13g2_inv_1 _04639_ (.VDD(VPWR),
    .Y(_01401_),
    .A(\i_exotiny._2034_[3] ),
    .VSS(VGND));
 sg13g2_inv_2 _04640_ (.Y(_01402_),
    .A(net3780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _04641_ (.Y(_01403_),
    .A(net3768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _04642_ (.Y(_01404_),
    .A(\i_exotiny._0369_[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04643_ (.VDD(VPWR),
    .Y(_01405_),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_2 _04644_ (.Y(_01406_),
    .A(net2997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04645_ (.VDD(VPWR),
    .Y(_01407_),
    .A(net3589),
    .VSS(VGND));
 sg13g2_inv_1 _04646_ (.VDD(VPWR),
    .Y(_01408_),
    .A(net1967),
    .VSS(VGND));
 sg13g2_inv_1 _04647_ (.VDD(VPWR),
    .Y(_01409_),
    .A(net1935),
    .VSS(VGND));
 sg13g2_inv_1 _04648_ (.VDD(VPWR),
    .Y(_01410_),
    .A(net1968),
    .VSS(VGND));
 sg13g2_inv_1 _04649_ (.VDD(VPWR),
    .Y(_01411_),
    .A(\i_exotiny.i_wb_spi.dat_rx_r[8] ),
    .VSS(VGND));
 sg13g2_inv_1 _04650_ (.VDD(VPWR),
    .Y(_01412_),
    .A(net2105),
    .VSS(VGND));
 sg13g2_inv_1 _04651_ (.VDD(VPWR),
    .Y(_01413_),
    .A(net1897),
    .VSS(VGND));
 sg13g2_inv_1 _04652_ (.VDD(VPWR),
    .Y(_01414_),
    .A(net1905),
    .VSS(VGND));
 sg13g2_inv_2 _04653_ (.Y(_01415_),
    .A(net3777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04654_ (.VDD(VPWR),
    .Y(_01416_),
    .A(net1951),
    .VSS(VGND));
 sg13g2_inv_2 _04655_ (.Y(_01417_),
    .A(\i_exotiny.i_wb_spi.dat_rx_r[17] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04656_ (.VDD(VPWR),
    .Y(_01418_),
    .A(net2),
    .VSS(VGND));
 sg13g2_inv_1 _04657_ (.VDD(VPWR),
    .Y(_01419_),
    .A(net4),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _04659_ (.A(net1252),
    .B_N(net1250),
    .Y(_01420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _04660_ (.A(net1247),
    .B_N(_01420_),
    .Y(_01421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _04661_ (.Y(_01422_),
    .B(_01420_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1247));
 sg13g2_nor2_2 _04662_ (.A(net1242),
    .B(net1247),
    .Y(_01423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04663_ (.A(_01420_),
    .B(_01423_),
    .X(_01424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04664_ (.Y(_01425_),
    .A(_01420_),
    .B(_01423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04665_ (.A(net3692),
    .B(net3822),
    .C(net3670),
    .Y(_01426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _04666_ (.A(net1252),
    .B(net1253),
    .Y(_01427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04667_ (.A(net1250),
    .B(net1252),
    .C(net1253),
    .Y(_01428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04668_ (.A(net1249),
    .B(net1247),
    .C(net1243),
    .Y(_01429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04669_ (.A(_01428_),
    .B(_01429_),
    .X(_01430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04670_ (.A(net1242),
    .B(net1245),
    .C(net1247),
    .Y(_01431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04671_ (.A(net1248),
    .B(net1254),
    .Y(_01432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _04672_ (.A(net1248),
    .B(net1250),
    .C(net1252),
    .Y(_01433_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1253));
 sg13g2_a22oi_1 _04673_ (.Y(_01434_),
    .B1(_01431_),
    .B2(_01433_),
    .A2(_01429_),
    .A1(_01428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _04674_ (.A2(_01433_),
    .A1(_01431_),
    .B1(_01430_),
    .X(_01435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04675_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0315_[8] ),
    .A2(net1201),
    .Y(_01436_),
    .B1(_01430_));
 sg13g2_nor2_2 _04676_ (.A(\i_exotiny._0327_[0] ),
    .B(net1234),
    .Y(_01437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04677_ (.Y(_01438_),
    .B1(_01435_),
    .B2(net3790),
    .A2(_01426_),
    .A1(_01424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04678_ (.A(net3523),
    .B(net3677),
    .C(net1984),
    .Y(_01439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _04679_ (.B(_01439_),
    .A(net3827),
    .X(_01440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04680_ (.Y(_01441_),
    .A(net1266),
    .B(_01440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04681_ (.B1(_01441_),
    .VDD(VPWR),
    .Y(\i_exotiny._1489_[3] ),
    .VSS(VGND),
    .A1(net1266),
    .A2(_01438_));
 sg13g2_nand2_1 _04682_ (.Y(_01442_),
    .A(net3832),
    .B(net3824),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04683_ (.B(net3832),
    .C(net3824),
    .A(net3834),
    .Y(_01443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _04684_ (.Y(\i_exotiny._1265_ ),
    .A(_01443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04685_ (.B1(net1281),
    .VDD(VPWR),
    .Y(_01444_),
    .VSS(VGND),
    .A1(_01364_),
    .A2(net3241));
 sg13g2_nor2_1 _04686_ (.A(net1266),
    .B(\i_exotiny._0315_[6] ),
    .Y(_01445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04687_ (.Y(\i_exotiny._1489_[0] ),
    .B1(net1202),
    .B2(_01445_),
    .A2(net3523),
    .A1(net1266),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04688_ (.A(\i_exotiny._1489_[3] ),
    .B(\i_exotiny._1489_[0] ),
    .X(_01446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _04689_ (.A0(\i_exotiny._0315_[29] ),
    .A1(\i_exotiny._0314_[29] ),
    .S(net1271),
    .X(_01447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04690_ (.Y(_01448_),
    .A(net1270),
    .B(_01447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04691_ (.A(\i_exotiny._0315_[30] ),
    .B(net1278),
    .Y(_01449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _04692_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_01449_),
    .Y(_01450_),
    .A2(net1279),
    .A1(_01370_));
 sg13g2_a21o_2 _04693_ (.A2(net1279),
    .A1(_01370_),
    .B1(_01449_),
    .X(_01451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04694_ (.A(net3705),
    .B(net3841),
    .Y(_01452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04695_ (.B(net1187),
    .C(_01452_),
    .A(_01448_),
    .Y(_01453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04696_ (.A(net1270),
    .B(_01453_),
    .X(_01454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04697_ (.B1(_01446_),
    .VDD(VPWR),
    .Y(_01455_),
    .VSS(VGND),
    .A1(net1266),
    .A2(_01454_));
 sg13g2_nand2_1 _04698_ (.Y(_01456_),
    .A(net1248),
    .B(net1247),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04699_ (.A(net1251),
    .B(_01456_),
    .Y(_01457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04700_ (.A(net1251),
    .B(net1252),
    .C(_01456_),
    .Y(_01458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04701_ (.A(net1224),
    .B(_01458_),
    .X(_01459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _04702_ (.A2(_01458_),
    .A1(net1242),
    .B1(_01459_),
    .X(_01460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _04703_ (.A(net1253),
    .B_N(_01460_),
    .Y(_01461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04704_ (.Y(_01462_),
    .A(net1245),
    .B(net1243),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04705_ (.A(_01423_),
    .B(_01428_),
    .X(_01463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _04706_ (.X(_01464_),
    .A(net1249),
    .B(_01462_),
    .C(_01463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04707_ (.B(_01462_),
    .C(_01463_),
    .A(net1249),
    .Y(_01465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04708_ (.A(net1253),
    .B(_01457_),
    .X(_01466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04709_ (.Y(_01467_),
    .A(net1253),
    .B(_01457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04710_ (.Y(_01468_),
    .A(net1243),
    .B(_01421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04711_ (.A(net1254),
    .B(_01468_),
    .Y(_01469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04712_ (.A(\i_exotiny._0571_ ),
    .B(net1253),
    .C(_01468_),
    .Y(_01470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _04713_ (.A(_01461_),
    .B(_01464_),
    .C(_01466_),
    .D(_01470_),
    .Y(_01471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _04714_ (.A(\i_exotiny._0590_ ),
    .B(net1250),
    .C(net1252),
    .D(_01432_),
    .X(_01472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _04715_ (.B(net1251),
    .C(net1252),
    .A(\i_exotiny._0590_ ),
    .Y(_01473_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01432_));
 sg13g2_nor2_1 _04716_ (.A(net14),
    .B(_01473_),
    .Y(_01474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04717_ (.A(_01443_),
    .B(_01474_),
    .Y(_01475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04718_ (.VDD(VPWR),
    .Y(_01476_),
    .A(_01475_),
    .VSS(VGND));
 sg13g2_nand2_1 _04719_ (.Y(_01477_),
    .A(net3819),
    .B(_01475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _04720_ (.Y(_01478_),
    .A(_01477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04721_ (.A(net1174),
    .B(_01471_),
    .C(_01477_),
    .Y(_01479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04722_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1269),
    .A2(_01443_),
    .Y(_01480_),
    .B1(_01479_));
 sg13g2_a21oi_1 _04723_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01455_),
    .A2(_01480_),
    .Y(_00004_),
    .B1(net1197));
 sg13g2_nand3_1 _04724_ (.B(\i_exotiny._1265_ ),
    .C(_01464_),
    .A(net1268),
    .Y(_01481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04725_ (.B1(_01481_),
    .VDD(VPWR),
    .Y(_01482_),
    .VSS(VGND),
    .A1(_01380_),
    .A2(_01453_));
 sg13g2_a21oi_1 _04726_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01435_),
    .A2(_01478_),
    .Y(_01483_),
    .B1(_01482_));
 sg13g2_nor2_1 _04727_ (.A(net1196),
    .B(_01483_),
    .Y(_00003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04728_ (.A(\i_exotiny._1309_ ),
    .B(_01464_),
    .X(_01484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04729_ (.Y(_01485_),
    .A(net3754),
    .B(_01464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04730_ (.Y(_01486_),
    .A(net1230),
    .B(net1231),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _04731_ (.X(_01487_),
    .A(net1230),
    .B(net1231),
    .C(net3713),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04732_ (.B(net1231),
    .C(net3713),
    .A(net1230),
    .Y(_01488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _04733_ (.A0(\i_exotiny._0315_[28] ),
    .A1(\i_exotiny._0314_[28] ),
    .S(net1271),
    .X(_01489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _04734_ (.B(net1231),
    .C(net3713),
    .A(_01383_),
    .Y(_01490_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net1218));
 sg13g2_a21oi_1 _04735_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01488_),
    .A2(_01490_),
    .Y(_01491_),
    .B1(net1226));
 sg13g2_nand2_1 _04736_ (.Y(_01492_),
    .A(net3724),
    .B(_01491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _04737_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01493_),
    .B(_01486_),
    .A(\i_exotiny.i_wb_qspi_mem.cnt_r[2] ));
 sg13g2_nand3_1 _04738_ (.B(net3520),
    .C(_01493_),
    .A(net1283),
    .Y(_01494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04739_ (.B1(net3521),
    .VDD(VPWR),
    .Y(_00007_),
    .VSS(VGND),
    .A1(net1146),
    .A2(_01492_));
 sg13g2_a21oi_1 _04740_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1306_ ),
    .A2(_01476_),
    .Y(_01495_),
    .B1(net1893));
 sg13g2_nor2_1 _04741_ (.A(net1197),
    .B(net1894),
    .Y(_00002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _04742_ (.A(net1243),
    .B(_01422_),
    .Y(_01496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04743_ (.A(net1245),
    .B(_01421_),
    .X(_01497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04744_ (.Y(_01498_),
    .A(net1245),
    .B(_01421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04745_ (.A(net1254),
    .B(net1243),
    .C(_01498_),
    .Y(_01499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _04746_ (.B(net1224),
    .C(_01497_),
    .Y(_01500_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1254));
 sg13g2_nand4_1 _04747_ (.B(_01471_),
    .C(_01478_),
    .A(net1202),
    .Y(_01501_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01500_));
 sg13g2_nand3_1 _04748_ (.B(\i_exotiny._1265_ ),
    .C(_01465_),
    .A(net1268),
    .Y(_01502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04749_ (.A(net1279),
    .B(\i_exotiny._1623_ ),
    .X(_01503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04750_ (.Y(_01504_),
    .A(net1279),
    .B(net3705),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _04751_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net1273),
    .C1(net1196),
    .B1(net1212),
    .A1(net1201),
    .Y(_01505_),
    .A2(_01454_));
 sg13g2_nand3_1 _04752_ (.B(_01502_),
    .C(_01505_),
    .A(_01501_),
    .Y(_00001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _04753_ (.A2(_01488_),
    .A1(net3651),
    .B1(net1226),
    .X(_00006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04754_ (.A(net1174),
    .B(_01454_),
    .X(_01506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04755_ (.Y(_01507_),
    .A(net1174),
    .B(_01454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _04756_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01499_),
    .C1(net3694),
    .B1(_01478_),
    .A1(net1174),
    .Y(_01508_),
    .A2(_01454_));
 sg13g2_nor3_1 _04757_ (.A(net1196),
    .B(_01446_),
    .C(net3695),
    .Y(_00005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04758_ (.A(net1230),
    .B(_01384_),
    .C(\i_exotiny.i_wb_qspi_mem.cnt_r[2] ),
    .Y(_01509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _04759_ (.A2(_01509_),
    .A1(net1218),
    .B1(_01487_),
    .X(_01510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _04760_ (.VDD(VPWR),
    .Y(_01511_),
    .A(_01510_),
    .VSS(VGND));
 sg13g2_and2_1 _04761_ (.A(net1265),
    .B(_01510_),
    .X(_01512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04762_ (.Y(_01513_),
    .A(net1265),
    .B(_01510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04763_ (.A(net1272),
    .B(\i_exotiny._0315_[31] ),
    .Y(_01514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _04764_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_01514_),
    .Y(_01515_),
    .A2(net1271),
    .A1(_01369_));
 sg13g2_nor2_1 _04765_ (.A(net1219),
    .B(net1181),
    .Y(_01516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _04766_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01517_),
    .B(net1181),
    .A(net1219));
 sg13g2_nor2_1 _04767_ (.A(net1270),
    .B(net1273),
    .Y(_01518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04768_ (.A(net1193),
    .B(net1169),
    .C(_01518_),
    .Y(_01519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04769_ (.A(net3830),
    .B(_01519_),
    .X(_01520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04770_ (.Y(_01521_),
    .A(net3830),
    .B(_01519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _04771_ (.Y(_01522_),
    .B(net3775),
    .A_N(net1218),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04772_ (.B1(_01513_),
    .VDD(VPWR),
    .Y(_01523_),
    .VSS(VGND),
    .A1(_01521_),
    .A2(_01522_));
 sg13g2_nand2_1 _04773_ (.Y(_01524_),
    .A(net1146),
    .B(_01513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04774_ (.A(_01523_),
    .B(_01524_),
    .X(_01525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04775_ (.Y(_01526_),
    .A(net1283),
    .B(_01525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _04776_ (.X(_01527_),
    .A(net3724),
    .B(_01488_),
    .C(_01490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04777_ (.A(_01525_),
    .B(_01527_),
    .Y(_01528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04778_ (.A(net1226),
    .B(_01528_),
    .Y(_00012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04779_ (.Y(_01529_),
    .A(net1224),
    .B(net1234),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04780_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1246),
    .A2(_01387_),
    .Y(_01530_),
    .B1(net1273));
 sg13g2_nor2b_1 _04781_ (.A(_01529_),
    .B_N(_01530_),
    .Y(_01531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04782_ (.A(net1246),
    .B(net1244),
    .Y(_01532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _04783_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01533_),
    .B(net1244),
    .A(net1246));
 sg13g2_a221oi_1 _04784_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01533_),
    .C1(net1273),
    .B1(_01437_),
    .A1(net1224),
    .Y(_01534_),
    .A2(net1234));
 sg13g2_xnor2_1 _04785_ (.Y(_01535_),
    .A(net1230),
    .B(_01534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04786_ (.A(net1273),
    .B(_01437_),
    .Y(_01536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04787_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1243),
    .A2(_01437_),
    .Y(_01537_),
    .B1(net1273));
 sg13g2_xor2_1 _04788_ (.B(_01537_),
    .A(net3713),
    .X(_01538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _04789_ (.Y(_01539_),
    .A(_01531_),
    .B(_01535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04790_ (.B(_01538_),
    .C(_01539_),
    .A(net1231),
    .Y(_01540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04791_ (.Y(_01541_),
    .A(net1283),
    .B(net1264),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04792_ (.B(net3702),
    .C(_01487_),
    .A(net1281),
    .Y(_01542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04793_ (.B1(_01542_),
    .VDD(VPWR),
    .Y(_00013_),
    .VSS(VGND),
    .A1(_01540_),
    .A2(_01541_));
 sg13g2_nand2_1 _04794_ (.Y(_01543_),
    .A(net1283),
    .B(net3702),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _04795_ (.B(net1230),
    .C(net1232),
    .A(net1283),
    .Y(_01544_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net3520));
 sg13g2_a21oi_1 _04796_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01543_),
    .A2(_01544_),
    .Y(_00011_),
    .B1(_01487_));
 sg13g2_nor2b_1 _04797_ (.A(_01519_),
    .B_N(\i_exotiny._1757_ ),
    .Y(_01545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04798_ (.B1(net1283),
    .VDD(VPWR),
    .Y(_01546_),
    .VSS(VGND),
    .A1(\i_exotiny._1623_ ),
    .A2(_01545_));
 sg13g2_nand3_1 _04799_ (.B(net3651),
    .C(_01487_),
    .A(net1282),
    .Y(_01547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04800_ (.Y(_00010_),
    .A(_01546_),
    .B(net3652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04801_ (.Y(_01548_),
    .A(net1270),
    .B(net1181),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _04802_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01549_),
    .B(_01548_),
    .A(\i_exotiny._3871_ ));
 sg13g2_inv_2 _04803_ (.Y(_00026_),
    .A(net1144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04804_ (.A(\i_exotiny._0315_[2] ),
    .B(_01549_),
    .Y(_01550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _04805_ (.Y(_01551_),
    .B(net1127),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1233));
 sg13g2_nor4_2 _04806_ (.A(net3789),
    .B(net1234),
    .C(_01465_),
    .Y(\i_exotiny._2160_ ),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01551_));
 sg13g2_nand2b_1 _04807_ (.Y(_01552_),
    .B(_01540_),
    .A_N(_01541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04808_ (.B1(_01552_),
    .VDD(VPWR),
    .Y(_00009_),
    .VSS(VGND),
    .A1(_01485_),
    .A2(_01492_));
 sg13g2_nor2_2 _04809_ (.A(_01485_),
    .B(_01521_),
    .Y(_01553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _04810_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01522_),
    .C1(_01553_),
    .B1(_01520_),
    .A1(net1265),
    .Y(_01554_),
    .A2(_01511_));
 sg13g2_nor2_1 _04811_ (.A(net1226),
    .B(_01554_),
    .Y(_00008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _04812_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01555_),
    .B(\i_exotiny._1757_ ),
    .A(\i_exotiny._1623_ ));
 sg13g2_a21oi_1 _04813_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1226),
    .A2(\i_exotiny._1793_ ),
    .Y(_01556_),
    .B1(_01555_));
 sg13g2_o21ai_1 _04814_ (.B1(_01556_),
    .VDD(VPWR),
    .Y(\i_exotiny._5416_$func$/home/user/heichips25-fazyrv-exotiny/build/exotiny_preproc.v:7385$12.$result [0]),
    .VSS(VGND),
    .A1(\i_exotiny._1793_ ),
    .A2(net1218));
 sg13g2_nor2_1 _04815_ (.A(\i_exotiny._1725_ ),
    .B(net1264),
    .Y(_01557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04816_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1281),
    .A2(\i_exotiny._1793_ ),
    .Y(_01558_),
    .B1(net1265));
 sg13g2_nand2_2 _04817_ (.Y(net19),
    .A(_01557_),
    .B(_01558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04818_ (.Y(_01559_),
    .A(net1265),
    .B(net1218),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04819_ (.Y(net22),
    .A(_01557_),
    .B(_01559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _04820_ (.A(net1852),
    .B(net1845),
    .C(net1856),
    .D(net1843),
    .Y(_01560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _04821_ (.A(net1867),
    .B(net1868),
    .C(net1865),
    .D(net1839),
    .Y(_01561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _04822_ (.A(\i_exotiny.i_wb_spi.state_r[24] ),
    .B(\i_exotiny.i_wb_spi.state_r[27] ),
    .C(\i_exotiny.i_wb_spi.state_r[26] ),
    .D(\i_exotiny.i_wb_spi.state_r[29] ),
    .X(_01562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _04823_ (.A(net1866),
    .B(net1854),
    .C(net1864),
    .D(_01562_),
    .Y(_01563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04824_ (.B(_01561_),
    .C(_01563_),
    .A(_01560_),
    .Y(_01564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _04825_ (.A(net1849),
    .B(net1841),
    .C(net1835),
    .D(net1859),
    .X(_01565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _04826_ (.A(net1846),
    .B(net1858),
    .C(net1853),
    .D(net1837),
    .Y(_01566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _04827_ (.A(net1869),
    .B(net1857),
    .C(net1855),
    .D(net1847),
    .Y(_01567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _04828_ (.A(net1863),
    .B(net1851),
    .C(net1861),
    .D(net1848),
    .Y(_01568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04829_ (.B(_01567_),
    .C(_01568_),
    .A(_01566_),
    .Y(_01569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04830_ (.A(_01564_),
    .B(_01565_),
    .C(_01569_),
    .Y(_01570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04831_ (.Y(_01571_),
    .A(net3640),
    .B(_01570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04832_ (.A(net1840),
    .B(net3728),
    .C(net3814),
    .Y(_01572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _04833_ (.A(\i_exotiny.i_wb_spi.cnt_presc_r[3] ),
    .B_N(_01572_),
    .Y(_01573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _04834_ (.A(\i_exotiny.i_wb_spi.cnt_presc_r[4] ),
    .B_N(_01573_),
    .Y(_01574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _04835_ (.Y(_01575_),
    .B(_01574_),
    .A_N(\i_exotiny.i_wb_spi.cnt_presc_r[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04836_ (.A(\i_exotiny.i_wb_spi.cnt_presc_r[6] ),
    .B(_01575_),
    .Y(_01576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _04837_ (.A(_01571_),
    .B_N(_01576_),
    .Y(_01577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _04838_ (.A(net1187),
    .B(_01485_),
    .Y(_01578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04839_ (.Y(_01579_),
    .A(_01570_),
    .B(_01578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _04840_ (.A(net3634),
    .B(_01579_),
    .Y(_01580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04841_ (.A(net1111),
    .B(_01580_),
    .Y(_01581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04842_ (.A(_01379_),
    .B(_01570_),
    .X(_01582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04843_ (.A(_01578_),
    .B(net1118),
    .X(_01583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04844_ (.A(net1111),
    .B(_01583_),
    .Y(_01584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04845_ (.A(net1840),
    .B(net1111),
    .C(_01583_),
    .Y(\i_exotiny._1902_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _04846_ (.B(net3728),
    .A(net1840),
    .X(_01585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04847_ (.A(net1111),
    .B(_01583_),
    .C(_01585_),
    .Y(\i_exotiny._1902_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04848_ (.B1(net3814),
    .VDD(VPWR),
    .Y(_01586_),
    .VSS(VGND),
    .A1(net1840),
    .A2(net3728));
 sg13g2_nor2b_1 _04849_ (.A(_01572_),
    .B_N(_01586_),
    .Y(_01587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04850_ (.A(net1111),
    .B(_01583_),
    .C(_01587_),
    .Y(\i_exotiny._1902_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _04851_ (.Y(_01588_),
    .A(\i_exotiny.i_wb_spi.cnt_presc_r[3] ),
    .B(_01572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04852_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3551),
    .A2(_01570_),
    .Y(_01589_),
    .B1(net1072));
 sg13g2_a21oi_1 _04853_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1072),
    .A2(_01588_),
    .Y(\i_exotiny._1902_[3] ),
    .B1(_01589_));
 sg13g2_xnor2_1 _04854_ (.Y(_01590_),
    .A(\i_exotiny.i_wb_spi.cnt_presc_r[4] ),
    .B(_01573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04855_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3618),
    .A2(_01570_),
    .Y(_01591_),
    .B1(net1072));
 sg13g2_a21oi_1 _04856_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1072),
    .A2(_01590_),
    .Y(\i_exotiny._1902_[4] ),
    .B1(_01591_));
 sg13g2_xnor2_1 _04857_ (.Y(_01592_),
    .A(\i_exotiny.i_wb_spi.cnt_presc_r[5] ),
    .B(_01574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04858_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3561),
    .A2(_01570_),
    .Y(_01593_),
    .B1(net1072));
 sg13g2_a21oi_1 _04859_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1072),
    .A2(_01592_),
    .Y(\i_exotiny._1902_[5] ),
    .B1(_01593_));
 sg13g2_and2_1 _04860_ (.A(_01571_),
    .B(_01576_),
    .X(_01594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04861_ (.Y(_01595_),
    .B1(_01579_),
    .B2(_01594_),
    .A2(_01575_),
    .A1(\i_exotiny.i_wb_spi.cnt_presc_r[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04862_ (.B1(net3430),
    .VDD(VPWR),
    .Y(_01596_),
    .VSS(VGND),
    .A1(net1111),
    .A2(_01583_));
 sg13g2_o21ai_1 _04863_ (.B1(_01596_),
    .VDD(VPWR),
    .Y(\i_exotiny._1902_[6] ),
    .VSS(VGND),
    .A1(_01580_),
    .A2(_01595_));
 sg13g2_nand2_1 _04864_ (.Y(_01597_),
    .A(net1266),
    .B(_01446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _04865_ (.A(net1268),
    .B(\i_exotiny._1306_ ),
    .Y(_01598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04866_ (.A(net1270),
    .B(net1267),
    .Y(_01599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _04867_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01599_),
    .C1(_01454_),
    .B1(_01598_),
    .A1(net1269),
    .Y(_01600_),
    .A2(\i_exotiny._1265_ ));
 sg13g2_nand3_1 _04868_ (.B(_01597_),
    .C(_01600_),
    .A(_01477_),
    .Y(\i_exotiny._1266_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04869_ (.A(net1271),
    .B(net1267),
    .C(net1268),
    .Y(_01601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _04870_ (.A(net1271),
    .B(net1266),
    .C(net1268),
    .X(_01602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04871_ (.B(_01381_),
    .C(_01427_),
    .A(net1248),
    .Y(_01603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04872_ (.B(net1250),
    .C(_01427_),
    .A(net1248),
    .Y(_01604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04873_ (.A(net1242),
    .B(_01604_),
    .Y(_01605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _04874_ (.A2(_01605_),
    .A1(net1247),
    .B1(_01499_),
    .X(_01606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _04875_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_01466_),
    .Y(_01607_),
    .A2(_01606_),
    .A1(_01601_));
 sg13g2_a21o_1 _04876_ (.A2(_01606_),
    .A1(_01601_),
    .B1(_01466_),
    .X(_01608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04877_ (.B1(_01466_),
    .VDD(VPWR),
    .Y(_01609_),
    .VSS(VGND),
    .A1(net1252),
    .A2(_01602_));
 sg13g2_nand2_1 _04878_ (.Y(_01610_),
    .A(net1254),
    .B(_01421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04879_ (.Y(_01611_),
    .B1(_01460_),
    .B2(_01602_),
    .A2(_01421_),
    .A1(net1254),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04880_ (.Y(_01612_),
    .A(_01609_),
    .B(_01611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _04881_ (.Y(_01613_),
    .B(net1258),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1260));
 sg13g2_or3_1 _04882_ (.A(\i_exotiny._0077_[2] ),
    .B(\i_exotiny._0077_[3] ),
    .C(net1223),
    .X(_01614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _04883_ (.A(_01613_),
    .B(_01614_),
    .Y(_01615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _04884_ (.Y(_01616_),
    .B(\i_exotiny._0077_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\i_exotiny._0077_[2] ));
 sg13g2_nand2_2 _04885_ (.Y(_01617_),
    .A(net1258),
    .B(net1260),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04886_ (.A(net1222),
    .B(_01616_),
    .C(_01617_),
    .Y(_01618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _04887_ (.A(\i_exotiny._0077_[2] ),
    .B(\i_exotiny._0077_[3] ),
    .C(net1255),
    .Y(_01619_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01613_));
 sg13g2_nand2b_2 _04888_ (.Y(_01620_),
    .B(net1260),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1259));
 sg13g2_nor3_2 _04889_ (.A(net1256),
    .B(_01616_),
    .C(_01620_),
    .Y(_01621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _04890_ (.A(\i_exotiny._0077_[2] ),
    .B(\i_exotiny._0077_[3] ),
    .C(net1256),
    .Y(_01622_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01620_));
 sg13g2_nand2b_2 _04891_ (.Y(_01623_),
    .B(\i_exotiny._0077_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\i_exotiny._0077_[3] ));
 sg13g2_nor3_2 _04892_ (.A(net1256),
    .B(_01613_),
    .C(_01623_),
    .Y(_01624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04893_ (.A(net1223),
    .B(_01613_),
    .C(_01616_),
    .Y(_01625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04894_ (.A(net1256),
    .B(_01616_),
    .C(_01617_),
    .Y(_01626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _04895_ (.A(net1258),
    .B(net1260),
    .C(net1222),
    .Y(_01627_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01616_));
 sg13g2_nor4_2 _04896_ (.A(\i_exotiny._0077_[2] ),
    .B(\i_exotiny._0077_[3] ),
    .C(net1257),
    .Y(_01628_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01617_));
 sg13g2_nand2_1 _04897_ (.Y(_01629_),
    .A(\i_exotiny._0037_[3] ),
    .B(_01628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04898_ (.A(net1256),
    .B(_01617_),
    .C(_01623_),
    .Y(_01630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04899_ (.A(net1222),
    .B(_01617_),
    .C(_01623_),
    .Y(_01631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _04900_ (.A(_01614_),
    .B(_01617_),
    .Y(_01632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04901_ (.Y(_01633_),
    .B1(_01632_),
    .B2(\i_exotiny._0022_[3] ),
    .A2(_01631_),
    .A1(\i_exotiny._0027_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04902_ (.A(net1255),
    .B(_01613_),
    .C(_01616_),
    .Y(_01634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04903_ (.Y(_01635_),
    .A(\i_exotiny._0013_[3] ),
    .B(_01634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04904_ (.A(net1258),
    .B(net1260),
    .C(_01614_),
    .Y(_01636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _04905_ (.A(net1258),
    .B(net1260),
    .C(net1222),
    .Y(_01637_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01623_));
 sg13g2_nor3_2 _04906_ (.A(net1222),
    .B(_01616_),
    .C(_01620_),
    .Y(_01638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04907_ (.Y(_01639_),
    .B1(_01638_),
    .B2(\i_exotiny._0029_[3] ),
    .A2(_01637_),
    .A1(\i_exotiny._0024_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04908_ (.Y(_01640_),
    .A(\i_exotiny._0077_[2] ),
    .B(\i_exotiny._0077_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04909_ (.A(net1222),
    .B(_01613_),
    .C(_01640_),
    .Y(_01641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _04910_ (.A(net1258),
    .B(net1261),
    .C(net1256),
    .Y(_01642_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01640_));
 sg13g2_nor2_2 _04911_ (.A(_01617_),
    .B(_01640_),
    .Y(_01643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _04912_ (.Y(_01644_),
    .A(net1256),
    .B(_01643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04913_ (.A(net1222),
    .B(_01620_),
    .C(_01623_),
    .Y(_01645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04914_ (.A(net1255),
    .B(_01613_),
    .C(_01640_),
    .Y(_01646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _04915_ (.A(net1259),
    .B(net1261),
    .C(net1223),
    .Y(_01647_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01640_));
 sg13g2_nor3_2 _04916_ (.A(net1222),
    .B(_01620_),
    .C(_01640_),
    .Y(_01648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _04917_ (.A(net1258),
    .B(net1260),
    .C(net1255),
    .Y(_01649_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01616_));
 sg13g2_nor3_2 _04918_ (.A(net1255),
    .B(_01620_),
    .C(_01640_),
    .Y(_01650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04919_ (.A(net1256),
    .B(_01620_),
    .C(_01623_),
    .Y(_01651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04920_ (.A(net1255),
    .B(_01617_),
    .C(_01640_),
    .Y(_01652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _04921_ (.A(net1258),
    .B(net1260),
    .C(net1255),
    .Y(_01653_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01623_));
 sg13g2_nor2_2 _04922_ (.A(_01614_),
    .B(_01620_),
    .Y(_01654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _04923_ (.A(net1223),
    .B(_01613_),
    .C(_01623_),
    .Y(_01655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04924_ (.Y(_01656_),
    .B1(_01648_),
    .B2(\i_exotiny._0033_[3] ),
    .A2(_01646_),
    .A1(\i_exotiny._0017_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04925_ (.Y(_01657_),
    .B1(_01650_),
    .B2(\i_exotiny._0016_[3] ),
    .A2(_01625_),
    .A1(\i_exotiny._0030_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04926_ (.Y(_01658_),
    .B1(_01652_),
    .B2(\i_exotiny._0018_[3] ),
    .A2(_01649_),
    .A1(\i_exotiny._0042_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _04927_ (.B(_01639_),
    .C(_01656_),
    .A(_01633_),
    .Y(_01659_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01658_));
 sg13g2_a22oi_1 _04928_ (.Y(_01660_),
    .B1(_01654_),
    .B2(\i_exotiny._0020_[3] ),
    .A2(_01653_),
    .A1(\i_exotiny._0038_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04929_ (.Y(_01661_),
    .B1(_01636_),
    .B2(\i_exotiny._0019_[3] ),
    .A2(_01627_),
    .A1(\i_exotiny._0028_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _04930_ (.B(_01657_),
    .C(_01660_),
    .A(_01635_),
    .Y(_01662_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01661_));
 sg13g2_a22oi_1 _04931_ (.Y(_01663_),
    .B1(_01624_),
    .B2(\i_exotiny._0040_[3] ),
    .A2(_01619_),
    .A1(\i_exotiny._0034_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04932_ (.Y(_01664_),
    .B1(_01630_),
    .B2(\i_exotiny._0041_[3] ),
    .A2(_01626_),
    .A1(\i_exotiny._0014_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04933_ (.Y(_01665_),
    .A(_01663_),
    .B(_01664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _04934_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0025_[3] ),
    .C1(_01665_),
    .B1(_01645_),
    .A1(\i_exotiny._0023_[3] ),
    .Y(_01666_),
    .A2(_01622_));
 sg13g2_a22oi_1 _04935_ (.Y(_01667_),
    .B1(_01641_),
    .B2(\i_exotiny._0035_[3] ),
    .A2(_01615_),
    .A1(\i_exotiny._0021_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04936_ (.Y(_01668_),
    .B1(_01655_),
    .B2(\i_exotiny._0026_[3] ),
    .A2(_01642_),
    .A1(\i_exotiny._0015_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04937_ (.Y(_01669_),
    .B1(_01621_),
    .B2(\i_exotiny._0043_[3] ),
    .A2(_01618_),
    .A1(\i_exotiny._0031_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04938_ (.B(_01668_),
    .C(_01669_),
    .A(_01667_),
    .Y(_01670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _04939_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0039_[3] ),
    .C1(_01670_),
    .B1(_01651_),
    .A1(\i_exotiny._0032_[3] ),
    .Y(_01671_),
    .A2(_01647_));
 sg13g2_nand4_1 _04940_ (.B(_01644_),
    .C(_01666_),
    .A(_01629_),
    .Y(_01672_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01671_));
 sg13g2_nor3_2 _04941_ (.A(_01659_),
    .B(_01662_),
    .C(_01672_),
    .Y(_01673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04942_ (.A(\i_exotiny._0036_[3] ),
    .B(_01644_),
    .Y(_01674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _04943_ (.A(_01612_),
    .B(_01673_),
    .C(_01674_),
    .Y(_01675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _04944_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_01675_),
    .Y(_01676_),
    .A2(_01612_),
    .A1(\i_exotiny._0314_[3] ));
 sg13g2_and2_1 _04945_ (.A(net1109),
    .B(_01676_),
    .X(_01677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04946_ (.A(net1245),
    .B(_01422_),
    .Y(_01678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04947_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1245),
    .A2(net1224),
    .Y(_01679_),
    .B1(net1248));
 sg13g2_nor3_1 _04948_ (.A(net1242),
    .B(_01533_),
    .C(_01604_),
    .Y(_01680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04949_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1242),
    .A2(net1184),
    .Y(_01681_),
    .B1(_01466_));
 sg13g2_a22oi_1 _04950_ (.Y(_01682_),
    .B1(_01680_),
    .B2(net1247),
    .A2(_01679_),
    .A1(_01421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04951_ (.Y(_01683_),
    .A(_01427_),
    .B(_01429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _04952_ (.Y(_01684_),
    .B1(_01462_),
    .B2(_01463_),
    .A2(_01429_),
    .A1(_01427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _04953_ (.Y(_01685_),
    .B(_01601_),
    .A_N(_01684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _04954_ (.B(_01681_),
    .C(_01682_),
    .A(_01611_),
    .Y(_01686_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01685_));
 sg13g2_mux2_1 _04955_ (.A0(_01532_),
    .A1(\i_exotiny._0315_[7] ),
    .S(net1201),
    .X(_01687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _04956_ (.Y(_01688_),
    .A(_01425_),
    .B(_01687_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04957_ (.Y(_01689_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ),
    .B(_01688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04958_ (.B(_01420_),
    .C(_01423_),
    .A(\i_exotiny._0315_[6] ),
    .Y(_01690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _04959_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01433_),
    .C1(_01386_),
    .B1(_01431_),
    .A1(_01428_),
    .Y(_01691_),
    .A2(_01429_));
 sg13g2_o21ai_1 _04960_ (.B1(_01690_),
    .VDD(VPWR),
    .Y(_01692_),
    .VSS(VGND),
    .A1(_01424_),
    .A2(_01691_));
 sg13g2_nand2_1 _04961_ (.Y(_01693_),
    .A(_01363_),
    .B(_01692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04962_ (.B1(_01693_),
    .VDD(VPWR),
    .Y(_01694_),
    .VSS(VGND),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ),
    .A2(_01688_));
 sg13g2_xor2_1 _04963_ (.B(_01688_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ),
    .X(_01695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _04964_ (.Y(_01696_),
    .A(_01424_),
    .B(_01436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _04965_ (.Y(_01697_),
    .B(_01362_),
    .A_N(_01696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _04966_ (.Y(_01698_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2] ),
    .B(_01696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04967_ (.A(_01363_),
    .B(_01692_),
    .Y(_01699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04968_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2] ),
    .A2(_01696_),
    .Y(_01700_),
    .B1(_01699_));
 sg13g2_nand4_1 _04969_ (.B(_01695_),
    .C(_01697_),
    .A(_01693_),
    .Y(_01701_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01700_));
 sg13g2_inv_1 _04970_ (.VDD(VPWR),
    .Y(_01702_),
    .A(_01701_),
    .VSS(VGND));
 sg13g2_nand3_1 _04971_ (.B(_01420_),
    .C(_01423_),
    .A(\i_exotiny._0315_[4] ),
    .Y(_01703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _04972_ (.Y(_01704_),
    .A(\i_exotiny._0315_[5] ),
    .B(_01703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _04973_ (.Y(_01705_),
    .A(_01393_),
    .B(_01703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _04974_ (.A(net1174),
    .B(_01705_),
    .Y(_01706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _04975_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01433_),
    .C1(_01391_),
    .B1(_01431_),
    .A1(_01428_),
    .Y(_01707_),
    .A2(_01429_));
 sg13g2_a221oi_1 _04976_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01433_),
    .C1(_01393_),
    .B1(_01431_),
    .A1(_01428_),
    .Y(_01708_),
    .A2(_01429_));
 sg13g2_nor2_1 _04977_ (.A(net1180),
    .B(_01708_),
    .Y(_01709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _04978_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01710_),
    .B(_01708_),
    .A(net1180));
 sg13g2_a21oi_1 _04979_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01424_),
    .A2(_01709_),
    .Y(_01711_),
    .B1(_01388_));
 sg13g2_o21ai_1 _04980_ (.B1(net1268),
    .VDD(VPWR),
    .Y(_01712_),
    .VSS(VGND),
    .A1(_01425_),
    .A2(_01710_));
 sg13g2_mux4_1 _04981_ (.S0(_01706_),
    .A0(\i_exotiny._6090_[0] ),
    .A1(\i_exotiny._6090_[2] ),
    .A2(\i_exotiny._6090_[1] ),
    .A3(\i_exotiny._6090_[3] ),
    .S1(net1180),
    .X(_01713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04982_ (.A(_01712_),
    .B(_01713_),
    .Y(_01714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04983_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01361_),
    .A2(_01712_),
    .Y(_01715_),
    .B1(_01714_));
 sg13g2_nor2_1 _04984_ (.A(net1242),
    .B(net1250),
    .Y(_01716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04985_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1250),
    .A2(\i_exotiny._0550_ ),
    .Y(_01717_),
    .B1(_01716_));
 sg13g2_mux4_1 _04986_ (.S0(net1180),
    .A0(\i_exotiny._6090_[2] ),
    .A1(\i_exotiny._6090_[3] ),
    .A2(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data [0]),
    .A3(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data [0]),
    .S1(_01706_),
    .X(_01718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04987_ (.A(_01712_),
    .B(_01718_),
    .Y(_01719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _04988_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01365_),
    .A2(_01712_),
    .Y(_01720_),
    .B1(_01719_));
 sg13g2_mux4_1 _04989_ (.S0(_01393_),
    .A0(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data [0]),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data [0]),
    .A2(_01713_),
    .A3(_01718_),
    .S1(_01711_),
    .X(_01721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _04990_ (.B(_01721_),
    .C(_01707_),
    .Y(_01722_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_01717_));
 sg13g2_mux2_1 _04991_ (.A0(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data [0]),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data [0]),
    .S(net1180),
    .X(_01723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _04992_ (.A0(\i_exotiny._6090_[3] ),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data [0]),
    .S(net1180),
    .X(_01724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04993_ (.B(_01704_),
    .C(_01723_),
    .A(net1201),
    .Y(_01725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _04994_ (.B1(_01724_),
    .VDD(VPWR),
    .Y(_01726_),
    .VSS(VGND),
    .A1(net1174),
    .A2(_01705_));
 sg13g2_nand3_1 _04995_ (.B(_01725_),
    .C(_01726_),
    .A(_01711_),
    .Y(_01727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _04996_ (.Y(_01728_),
    .B(_01712_),
    .A_N(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _04997_ (.A(_01727_),
    .B(_01728_),
    .X(_01729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _04998_ (.B(_01727_),
    .C(_01728_),
    .A(_01709_),
    .Y(_01730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _04999_ (.A(_01392_),
    .B(net1180),
    .Y(_01731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05000_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._6090_[2] ),
    .C1(_01731_),
    .B1(net1180),
    .A1(net1201),
    .Y(_01732_),
    .A2(_01704_));
 sg13g2_nor3_1 _05001_ (.A(net1174),
    .B(_01705_),
    .C(_01724_),
    .Y(_01733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05002_ (.B1(_01711_),
    .VDD(VPWR),
    .Y(_01734_),
    .VSS(VGND),
    .A1(_01732_),
    .A2(_01733_));
 sg13g2_nand2_1 _05003_ (.Y(_01735_),
    .A(_01366_),
    .B(_01712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05004_ (.A(_01734_),
    .B(_01735_),
    .X(_01736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05005_ (.B(_01708_),
    .C(_01734_),
    .A(_01391_),
    .Y(_01737_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01735_));
 sg13g2_a21o_1 _05006_ (.A2(_01737_),
    .A1(_01730_),
    .B1(_01717_),
    .X(_01738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _05007_ (.A2(_01738_),
    .A1(_01722_),
    .B1(_01701_),
    .X(_01739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05008_ (.B(_01694_),
    .C(_01698_),
    .A(_01689_),
    .Y(_01740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05009_ (.B(_01701_),
    .C(_01740_),
    .A(_01697_),
    .Y(_01741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _05010_ (.Y(_01742_),
    .A(_01424_),
    .B(_01741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05011_ (.B(_01739_),
    .C(_01742_),
    .A(_01371_),
    .Y(_01743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _05012_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01744_),
    .B(_01742_),
    .A(_01729_));
 sg13g2_a21oi_1 _05013_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01743_),
    .A2(_01744_),
    .Y(_01745_),
    .B1(_01702_));
 sg13g2_nand2_1 _05014_ (.Y(_01746_),
    .A(_01425_),
    .B(_01710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05015_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01371_),
    .A2(_01739_),
    .Y(_01747_),
    .B1(_01746_));
 sg13g2_a21o_1 _05016_ (.A2(_01746_),
    .A1(_01729_),
    .B1(_01701_),
    .X(_01748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05017_ (.B1(_01385_),
    .VDD(VPWR),
    .Y(_01749_),
    .VSS(VGND),
    .A1(_01747_),
    .A2(_01748_));
 sg13g2_o21ai_1 _05018_ (.B1(_01602_),
    .VDD(VPWR),
    .Y(_01750_),
    .VSS(VGND),
    .A1(net1174),
    .A2(_01499_));
 sg13g2_a21oi_1 _05019_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1267),
    .A2(\i_exotiny._6090_[3] ),
    .Y(_01751_),
    .B1(_01750_));
 sg13g2_o21ai_1 _05020_ (.B1(_01751_),
    .VDD(VPWR),
    .Y(_01752_),
    .VSS(VGND),
    .A1(_01745_),
    .A2(_01749_));
 sg13g2_nand2_2 _05021_ (.Y(_01753_),
    .A(net1238),
    .B(net1240),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _05022_ (.Y(_01754_),
    .A(\i_exotiny._0079_[2] ),
    .B(\i_exotiny._0079_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _05023_ (.A(net1221),
    .B(_01753_),
    .C(_01754_),
    .X(_01755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _05024_ (.Y(_01756_),
    .B(net1238),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1240));
 sg13g2_nand2b_2 _05025_ (.Y(_01757_),
    .B(\i_exotiny._0079_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\i_exotiny._0079_[3] ));
 sg13g2_nor3_2 _05026_ (.A(net1235),
    .B(_01756_),
    .C(_01757_),
    .Y(_01758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _05027_ (.Y(_01759_),
    .B(\i_exotiny._0079_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\i_exotiny._0079_[2] ));
 sg13g2_nor3_2 _05028_ (.A(net1235),
    .B(_01753_),
    .C(_01759_),
    .Y(_01760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _05029_ (.A(net1238),
    .B(net1240),
    .C(net1237),
    .Y(_01761_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01754_));
 sg13g2_nand2b_2 _05030_ (.Y(_01762_),
    .B(net1240),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1238));
 sg13g2_nor3_2 _05031_ (.A(net1220),
    .B(_01759_),
    .C(_01762_),
    .Y(_01763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05032_ (.Y(_01764_),
    .A(\i_exotiny._0029_[3] ),
    .B(_01763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05033_ (.A(net1220),
    .B(_01753_),
    .C(_01757_),
    .Y(_01765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05034_ (.A(net1220),
    .B(_01756_),
    .C(_01759_),
    .Y(_01766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _05035_ (.A(net1239),
    .B(net1240),
    .C(net1220),
    .Y(_01767_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01754_));
 sg13g2_or3_1 _05036_ (.A(\i_exotiny._0079_[2] ),
    .B(\i_exotiny._0079_[3] ),
    .C(net1221),
    .X(_01768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _05037_ (.A(_01753_),
    .B(_01768_),
    .Y(_01769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05038_ (.A(net1221),
    .B(_01757_),
    .C(_01762_),
    .Y(_01770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05039_ (.A(net1235),
    .B(_01754_),
    .C(_01762_),
    .Y(_01771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05040_ (.A(net1220),
    .B(_01754_),
    .C(_01762_),
    .Y(_01772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05041_ (.A(net1238),
    .B(net1240),
    .C(_01768_),
    .Y(_01773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05042_ (.A(net1236),
    .B(_01753_),
    .C(_01754_),
    .Y(_01774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05043_ (.Y(_01775_),
    .A(\i_exotiny._0018_[3] ),
    .B(_01774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _05044_ (.A(_01756_),
    .B(_01768_),
    .Y(_01776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05045_ (.A(net1235),
    .B(_01756_),
    .C(_01759_),
    .Y(_01777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05046_ (.A(net1220),
    .B(_01754_),
    .C(_01756_),
    .Y(_01778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _05047_ (.A(_01762_),
    .B(_01768_),
    .Y(_01779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05048_ (.A(net1236),
    .B(_01753_),
    .C(_01757_),
    .Y(_01780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _05049_ (.A(net1238),
    .B(net1240),
    .C(net1220),
    .Y(_01781_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01759_));
 sg13g2_nor4_2 _05050_ (.A(\i_exotiny._0079_[2] ),
    .B(\i_exotiny._0079_[3] ),
    .C(net1235),
    .Y(_01782_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01753_));
 sg13g2_nor4_2 _05051_ (.A(\i_exotiny._0079_[2] ),
    .B(\i_exotiny._0079_[3] ),
    .C(net1235),
    .Y(_01783_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01762_));
 sg13g2_nor4_2 _05052_ (.A(net1238),
    .B(net1241),
    .C(net1235),
    .Y(_01784_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01759_));
 sg13g2_nor3_2 _05053_ (.A(net1236),
    .B(_01759_),
    .C(_01762_),
    .Y(_01785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05054_ (.A(net1236),
    .B(_01754_),
    .C(_01756_),
    .Y(_01786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05055_ (.A(net1221),
    .B(_01753_),
    .C(_01759_),
    .Y(_01787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05056_ (.A(net1236),
    .B(_01757_),
    .C(_01762_),
    .Y(_01788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _05057_ (.A(net1238),
    .B(net1240),
    .C(net1220),
    .Y(_01789_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01757_));
 sg13g2_nor4_2 _05058_ (.A(\i_exotiny._0079_[2] ),
    .B(\i_exotiny._0079_[3] ),
    .C(net1235),
    .Y(_01790_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01756_));
 sg13g2_nor3_2 _05059_ (.A(net1221),
    .B(_01756_),
    .C(_01757_),
    .Y(_01791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _05060_ (.A(net1239),
    .B(net1241),
    .C(net1237),
    .Y(_01792_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01757_));
 sg13g2_a22oi_1 _05061_ (.Y(_01793_),
    .B1(_01791_),
    .B2(\i_exotiny._0026_[3] ),
    .A2(_01785_),
    .A1(\i_exotiny._0043_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05062_ (.Y(_01794_),
    .B1(_01790_),
    .B2(\i_exotiny._0034_[3] ),
    .A2(_01780_),
    .A1(\i_exotiny._0041_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05063_ (.Y(_01795_),
    .B1(_01784_),
    .B2(\i_exotiny._0042_[3] ),
    .A2(_01770_),
    .A1(\i_exotiny._0025_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05064_ (.Y(_01796_),
    .B1(_01773_),
    .B2(\i_exotiny._0019_[3] ),
    .A2(_01761_),
    .A1(\i_exotiny._0015_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05065_ (.Y(_01797_),
    .B1(_01783_),
    .B2(\i_exotiny._0023_[3] ),
    .A2(_01782_),
    .A1(\i_exotiny._0037_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05066_ (.Y(_01798_),
    .B1(_01786_),
    .B2(\i_exotiny._0017_[3] ),
    .A2(_01758_),
    .A1(\i_exotiny._0040_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05067_ (.B(_01796_),
    .C(_01797_),
    .A(_01793_),
    .Y(_01799_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01798_));
 sg13g2_a22oi_1 _05068_ (.Y(_01800_),
    .B1(_01789_),
    .B2(\i_exotiny._0024_[3] ),
    .A2(_01765_),
    .A1(\i_exotiny._0027_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05069_ (.B(_01794_),
    .C(_01795_),
    .A(_01775_),
    .Y(_01801_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01800_));
 sg13g2_nor2_1 _05070_ (.A(_01799_),
    .B(_01801_),
    .Y(_01802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05071_ (.Y(_01803_),
    .B1(_01787_),
    .B2(\i_exotiny._0031_[3] ),
    .A2(_01776_),
    .A1(\i_exotiny._0021_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05072_ (.Y(_01804_),
    .B1(_01792_),
    .B2(\i_exotiny._0038_[3] ),
    .A2(_01771_),
    .A1(\i_exotiny._0016_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05073_ (.B(_01764_),
    .C(_01803_),
    .A(_01755_),
    .Y(_01805_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01804_));
 sg13g2_a221oi_1 _05074_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0028_[3] ),
    .C1(_01805_),
    .B1(_01781_),
    .A1(\i_exotiny._0032_[3] ),
    .Y(_01806_),
    .A2(_01767_));
 sg13g2_a22oi_1 _05075_ (.Y(_01807_),
    .B1(_01788_),
    .B2(\i_exotiny._0039_[3] ),
    .A2(_01769_),
    .A1(\i_exotiny._0022_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05076_ (.Y(_01808_),
    .B1(_01778_),
    .B2(\i_exotiny._0035_[3] ),
    .A2(_01772_),
    .A1(\i_exotiny._0033_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05077_ (.Y(_01809_),
    .B1(_01779_),
    .B2(\i_exotiny._0020_[3] ),
    .A2(_01766_),
    .A1(\i_exotiny._0030_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05078_ (.B(_01808_),
    .C(_01809_),
    .A(_01807_),
    .Y(_01810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05079_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0013_[3] ),
    .C1(_01810_),
    .B1(_01777_),
    .A1(\i_exotiny._0014_[3] ),
    .Y(_01811_),
    .A2(_01760_));
 sg13g2_nand3_1 _05080_ (.B(_01806_),
    .C(_01811_),
    .A(_01802_),
    .Y(_01812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05081_ (.B1(_01812_),
    .VDD(VPWR),
    .Y(_01813_),
    .VSS(VGND),
    .A1(\i_exotiny._0036_[3] ),
    .A2(_01755_));
 sg13g2_a21oi_1 _05082_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01750_),
    .A2(_01813_),
    .Y(_01814_),
    .B1(net1108));
 sg13g2_a221oi_1 _05083_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01814_),
    .C1(net1109),
    .B1(_01752_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ),
    .Y(_01815_),
    .A2(net1107));
 sg13g2_nor2_1 _05084_ (.A(_01677_),
    .B(_01815_),
    .Y(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _05085_ (.Y(_01816_),
    .B(_01467_),
    .A_N(_01430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05086_ (.A(net1243),
    .B(_01603_),
    .Y(_01817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _05087_ (.Y(_01818_),
    .B(net1224),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_01603_));
 sg13g2_a21oi_1 _05088_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01428_),
    .A2(_01431_),
    .Y(_01819_),
    .B1(_01816_));
 sg13g2_o21ai_1 _05089_ (.B1(_01819_),
    .VDD(VPWR),
    .Y(_01820_),
    .VSS(VGND),
    .A1(net1250),
    .A2(_01818_));
 sg13g2_nor2_1 _05090_ (.A(net1248),
    .B(_01610_),
    .Y(_01821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _05091_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01822_),
    .B(_01821_),
    .A(_01680_));
 sg13g2_nor3_1 _05092_ (.A(net1245),
    .B(net1254),
    .C(_01422_),
    .Y(_01823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _05093_ (.A(_01461_),
    .B(_01469_),
    .C(_01822_),
    .D(_01823_),
    .X(_01824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _05094_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_01824_),
    .Y(_01825_),
    .A2(_01820_),
    .A1(_01601_));
 sg13g2_a221oi_1 _05095_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01814_),
    .C1(net1110),
    .B1(_01752_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ),
    .Y(_01826_),
    .A2(net1108));
 sg13g2_and2_1 _05096_ (.A(_01607_),
    .B(_01676_),
    .X(_01827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05097_ (.A(_01826_),
    .B(_01827_),
    .Y(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _05098_ (.A(_01825_),
    .B(_01826_),
    .C(_01827_),
    .X(_01828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05099_ (.A(net1248),
    .B(_01823_),
    .X(_01829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05100_ (.A(\i_exotiny._0550_ ),
    .B(_01829_),
    .X(_01830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _05101_ (.Y(_01831_),
    .A(\i_exotiny._0550_ ),
    .B(_01829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _05102_ (.A(_01677_),
    .B(_01815_),
    .C(_01830_),
    .X(_01832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05103_ (.B1(_01830_),
    .VDD(VPWR),
    .Y(_01833_),
    .VSS(VGND),
    .A1(_01677_),
    .A2(_01815_));
 sg13g2_a21o_2 _05104_ (.A2(_01833_),
    .A1(_01832_),
    .B1(_01828_),
    .X(_01834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05105_ (.B(_01832_),
    .C(_01833_),
    .A(_01828_),
    .Y(_01835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05106_ (.A(_01834_),
    .B(_01835_),
    .X(_01836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05107_ (.Y(_01837_),
    .A(_01834_),
    .B(_01835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _05108_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01838_),
    .B(_01742_),
    .A(_01720_));
 sg13g2_a21oi_1 _05109_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01743_),
    .A2(_01838_),
    .Y(_01839_),
    .B1(_01702_));
 sg13g2_o21ai_1 _05110_ (.B1(_01708_),
    .VDD(VPWR),
    .Y(_01840_),
    .VSS(VGND),
    .A1(\i_exotiny._0315_[4] ),
    .A2(_01425_));
 sg13g2_a21oi_1 _05111_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01371_),
    .A2(_01739_),
    .Y(_01841_),
    .B1(_01840_));
 sg13g2_a21o_1 _05112_ (.A2(_01840_),
    .A1(_01720_),
    .B1(_01701_),
    .X(_01842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05113_ (.B1(_01385_),
    .VDD(VPWR),
    .Y(_01843_),
    .VSS(VGND),
    .A1(_01841_),
    .A2(_01842_));
 sg13g2_a21oi_1 _05114_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1267),
    .A2(\i_exotiny._6090_[2] ),
    .Y(_01844_),
    .B1(_01750_));
 sg13g2_o21ai_1 _05115_ (.B1(_01844_),
    .VDD(VPWR),
    .Y(_01845_),
    .VSS(VGND),
    .A1(_01839_),
    .A2(_01843_));
 sg13g2_nor2_1 _05116_ (.A(\i_exotiny._0036_[2] ),
    .B(_01755_),
    .Y(_01846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05117_ (.Y(_01847_),
    .A(\i_exotiny._0032_[2] ),
    .B(_01767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05118_ (.Y(_01848_),
    .B1(_01783_),
    .B2(\i_exotiny._0023_[2] ),
    .A2(_01776_),
    .A1(\i_exotiny._0021_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05119_ (.Y(_01849_),
    .A(\i_exotiny._0019_[2] ),
    .B(_01773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05120_ (.Y(_01850_),
    .B1(_01784_),
    .B2(\i_exotiny._0042_[2] ),
    .A2(_01769_),
    .A1(\i_exotiny._0022_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05121_ (.Y(_01851_),
    .B1(_01771_),
    .B2(\i_exotiny._0016_[2] ),
    .A2(_01763_),
    .A1(\i_exotiny._0029_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05122_ (.Y(_01852_),
    .B1(_01772_),
    .B2(\i_exotiny._0033_[2] ),
    .A2(_01760_),
    .A1(\i_exotiny._0014_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05123_ (.Y(_01853_),
    .B1(_01789_),
    .B2(\i_exotiny._0024_[2] ),
    .A2(_01765_),
    .A1(\i_exotiny._0027_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05124_ (.Y(_01854_),
    .B1(_01777_),
    .B2(\i_exotiny._0013_[2] ),
    .A2(_01761_),
    .A1(\i_exotiny._0015_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05125_ (.B(_01852_),
    .C(_01853_),
    .A(_01850_),
    .Y(_01855_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01854_));
 sg13g2_a22oi_1 _05126_ (.Y(_01856_),
    .B1(_01788_),
    .B2(\i_exotiny._0039_[2] ),
    .A2(_01758_),
    .A1(\i_exotiny._0040_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05127_ (.Y(_01857_),
    .B1(_01792_),
    .B2(\i_exotiny._0038_[2] ),
    .A2(_01774_),
    .A1(\i_exotiny._0018_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05128_ (.B(_01851_),
    .C(_01856_),
    .A(_01847_),
    .Y(_01858_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01857_));
 sg13g2_a22oi_1 _05129_ (.Y(_01859_),
    .B1(_01790_),
    .B2(\i_exotiny._0034_[2] ),
    .A2(_01770_),
    .A1(\i_exotiny._0025_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05130_ (.Y(_01860_),
    .A(_01848_),
    .B(_01859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05131_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0031_[2] ),
    .C1(_01860_),
    .B1(_01787_),
    .A1(\i_exotiny._0020_[2] ),
    .Y(_01861_),
    .A2(_01779_));
 sg13g2_a22oi_1 _05132_ (.Y(_01862_),
    .B1(_01780_),
    .B2(\i_exotiny._0041_[2] ),
    .A2(_01778_),
    .A1(\i_exotiny._0035_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05133_ (.Y(_01863_),
    .B1(_01786_),
    .B2(\i_exotiny._0017_[2] ),
    .A2(_01782_),
    .A1(\i_exotiny._0037_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05134_ (.Y(_01864_),
    .B1(_01791_),
    .B2(\i_exotiny._0026_[2] ),
    .A2(_01785_),
    .A1(\i_exotiny._0043_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05135_ (.B(_01863_),
    .C(_01864_),
    .A(_01862_),
    .Y(_01865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05136_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0028_[2] ),
    .C1(_01865_),
    .B1(_01781_),
    .A1(\i_exotiny._0030_[2] ),
    .Y(_01866_),
    .A2(_01766_));
 sg13g2_nand4_1 _05137_ (.B(_01849_),
    .C(_01861_),
    .A(_01755_),
    .Y(_01867_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01866_));
 sg13g2_nor3_2 _05138_ (.A(_01855_),
    .B(_01858_),
    .C(_01867_),
    .Y(_01868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _05139_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01869_),
    .B(_01868_),
    .A(_01846_));
 sg13g2_a21oi_1 _05140_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01750_),
    .A2(_01869_),
    .Y(_01870_),
    .B1(net1108));
 sg13g2_and2_1 _05141_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ),
    .B(net1108),
    .X(_01871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _05142_ (.A2(_01870_),
    .A1(_01845_),
    .B1(_01871_),
    .X(_01872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05143_ (.Y(_01873_),
    .B1(_01642_),
    .B2(\i_exotiny._0015_[2] ),
    .A2(_01630_),
    .A1(\i_exotiny._0041_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05144_ (.Y(_01874_),
    .B1(_01626_),
    .B2(\i_exotiny._0014_[2] ),
    .A2(_01622_),
    .A1(\i_exotiny._0023_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05145_ (.Y(_01875_),
    .B1(_01641_),
    .B2(\i_exotiny._0035_[2] ),
    .A2(_01634_),
    .A1(\i_exotiny._0013_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05146_ (.Y(_01876_),
    .B1(_01654_),
    .B2(\i_exotiny._0020_[2] ),
    .A2(_01627_),
    .A1(\i_exotiny._0028_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05147_ (.Y(_01877_),
    .B1(_01646_),
    .B2(\i_exotiny._0017_[2] ),
    .A2(_01632_),
    .A1(\i_exotiny._0022_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05148_ (.B(_01876_),
    .C(_01877_),
    .A(_01874_),
    .Y(_01878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05149_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0039_[2] ),
    .C1(_01878_),
    .B1(_01651_),
    .A1(\i_exotiny._0034_[2] ),
    .Y(_01879_),
    .A2(_01619_));
 sg13g2_a22oi_1 _05150_ (.Y(_01880_),
    .B1(_01638_),
    .B2(\i_exotiny._0029_[2] ),
    .A2(_01625_),
    .A1(\i_exotiny._0030_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05151_ (.Y(_01881_),
    .B1(_01628_),
    .B2(\i_exotiny._0037_[2] ),
    .A2(_01624_),
    .A1(\i_exotiny._0040_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05152_ (.Y(_01882_),
    .A(_01873_),
    .B(_01881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05153_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0043_[2] ),
    .A2(_01621_),
    .Y(_01883_),
    .B1(_01882_));
 sg13g2_o21ai_1 _05154_ (.B1(_01643_),
    .VDD(VPWR),
    .Y(_01884_),
    .VSS(VGND),
    .A1(net1255),
    .A2(\i_exotiny._0018_[2] ));
 sg13g2_a22oi_1 _05155_ (.Y(_01885_),
    .B1(_01649_),
    .B2(\i_exotiny._0042_[2] ),
    .A2(_01647_),
    .A1(\i_exotiny._0032_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05156_ (.Y(_01886_),
    .B1(_01655_),
    .B2(\i_exotiny._0026_[2] ),
    .A2(_01615_),
    .A1(\i_exotiny._0021_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05157_ (.B(_01884_),
    .C(_01885_),
    .A(_01875_),
    .Y(_01887_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01886_));
 sg13g2_a22oi_1 _05158_ (.Y(_01888_),
    .B1(_01648_),
    .B2(\i_exotiny._0033_[2] ),
    .A2(_01631_),
    .A1(\i_exotiny._0027_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05159_ (.Y(_01889_),
    .B1(_01653_),
    .B2(\i_exotiny._0038_[2] ),
    .A2(_01618_),
    .A1(\i_exotiny._0031_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05160_ (.Y(_01890_),
    .B1(_01645_),
    .B2(\i_exotiny._0025_[2] ),
    .A2(_01637_),
    .A1(\i_exotiny._0024_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05161_ (.Y(_01891_),
    .B1(_01650_),
    .B2(\i_exotiny._0016_[2] ),
    .A2(_01636_),
    .A1(\i_exotiny._0019_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05162_ (.B(_01889_),
    .C(_01890_),
    .A(_01888_),
    .Y(_01892_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01891_));
 sg13g2_nor2_1 _05163_ (.A(_01887_),
    .B(_01892_),
    .Y(_01893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05164_ (.B(_01880_),
    .C(_01883_),
    .A(_01879_),
    .Y(_01894_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01893_));
 sg13g2_nor2_1 _05165_ (.A(\i_exotiny._0036_[2] ),
    .B(_01644_),
    .Y(_01895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05166_ (.A(_01612_),
    .B(_01895_),
    .Y(_01896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05167_ (.Y(_01897_),
    .B1(_01894_),
    .B2(_01896_),
    .A2(_01612_),
    .A1(\i_exotiny._0314_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05168_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01870_),
    .C1(net1110),
    .B1(_01845_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ),
    .Y(_01898_),
    .A2(net1107));
 sg13g2_and2_1 _05169_ (.A(net1110),
    .B(_01897_),
    .X(_01899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05170_ (.A(_01898_),
    .B(_01899_),
    .Y(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _05171_ (.A(_01825_),
    .B(_01898_),
    .C(_01899_),
    .X(_01900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05172_ (.A(net1110),
    .B(_01897_),
    .Y(_01901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05173_ (.A(net1109),
    .B(_01897_),
    .X(_01902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05174_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01870_),
    .C1(net1109),
    .B1(_01845_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ),
    .Y(_01903_),
    .A2(net1107));
 sg13g2_nor2_1 _05175_ (.A(_01902_),
    .B(_01903_),
    .Y(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05176_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01607_),
    .C1(_01901_),
    .B1(_01872_),
    .A1(\i_exotiny._0550_ ),
    .Y(_01904_),
    .A2(_01829_));
 sg13g2_o21ai_1 _05177_ (.B1(_01831_),
    .VDD(VPWR),
    .Y(_01905_),
    .VSS(VGND),
    .A1(_01902_),
    .A2(_01903_));
 sg13g2_nor3_1 _05178_ (.A(_01831_),
    .B(_01902_),
    .C(_01903_),
    .Y(_01906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _05179_ (.A(_01831_),
    .B(_01902_),
    .C(_01903_),
    .X(_01907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05180_ (.B1(_01900_),
    .VDD(VPWR),
    .Y(_01908_),
    .VSS(VGND),
    .A1(_01904_),
    .A2(_01906_));
 sg13g2_nor3_1 _05181_ (.A(_01900_),
    .B(_01904_),
    .C(_01906_),
    .Y(_01909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _05182_ (.B(_01905_),
    .C(_01907_),
    .Y(_01910_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_01900_));
 sg13g2_and2_1 _05183_ (.A(_01908_),
    .B(_01910_),
    .X(_01911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05184_ (.Y(_01912_),
    .B1(_01908_),
    .B2(_01910_),
    .A2(_01835_),
    .A1(_01834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _05185_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01913_),
    .B(_01742_),
    .A(_01736_));
 sg13g2_a21oi_1 _05186_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01743_),
    .A2(_01913_),
    .Y(_01914_),
    .B1(_01702_));
 sg13g2_o21ai_1 _05187_ (.B1(_01708_),
    .VDD(VPWR),
    .Y(_01915_),
    .VSS(VGND),
    .A1(\i_exotiny._0315_[4] ),
    .A2(_01424_));
 sg13g2_a21oi_1 _05188_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01371_),
    .A2(_01739_),
    .Y(_01916_),
    .B1(_01915_));
 sg13g2_a21o_1 _05189_ (.A2(_01915_),
    .A1(_01736_),
    .B1(_01701_),
    .X(_01917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05190_ (.B1(_01385_),
    .VDD(VPWR),
    .Y(_01918_),
    .VSS(VGND),
    .A1(_01916_),
    .A2(_01917_));
 sg13g2_a21oi_1 _05191_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1267),
    .A2(\i_exotiny._6090_[1] ),
    .Y(_01919_),
    .B1(_01750_));
 sg13g2_o21ai_1 _05192_ (.B1(_01919_),
    .VDD(VPWR),
    .Y(_01920_),
    .VSS(VGND),
    .A1(_01914_),
    .A2(_01918_));
 sg13g2_nand2_1 _05193_ (.Y(_01921_),
    .A(\i_exotiny._0024_[1] ),
    .B(_01789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05194_ (.Y(_01922_),
    .B1(_01777_),
    .B2(\i_exotiny._0013_[1] ),
    .A2(_01770_),
    .A1(\i_exotiny._0025_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05195_ (.Y(_01923_),
    .B1(_01781_),
    .B2(\i_exotiny._0028_[1] ),
    .A2(_01766_),
    .A1(\i_exotiny._0030_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05196_ (.Y(_01924_),
    .A(\i_exotiny._0035_[1] ),
    .B(_01778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05197_ (.Y(_01925_),
    .B1(_01786_),
    .B2(\i_exotiny._0017_[1] ),
    .A2(_01769_),
    .A1(\i_exotiny._0022_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05198_ (.Y(_01926_),
    .B1(_01782_),
    .B2(\i_exotiny._0037_[1] ),
    .A2(_01763_),
    .A1(\i_exotiny._0029_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05199_ (.Y(_01927_),
    .B1(_01779_),
    .B2(\i_exotiny._0020_[1] ),
    .A2(_01773_),
    .A1(\i_exotiny._0019_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05200_ (.Y(_01928_),
    .B1(_01787_),
    .B2(\i_exotiny._0031_[1] ),
    .A2(_01776_),
    .A1(\i_exotiny._0021_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05201_ (.Y(_01929_),
    .B1(_01780_),
    .B2(\i_exotiny._0041_[1] ),
    .A2(_01761_),
    .A1(\i_exotiny._0015_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05202_ (.B(_01925_),
    .C(_01928_),
    .A(_01923_),
    .Y(_01930_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01929_));
 sg13g2_a22oi_1 _05203_ (.Y(_01931_),
    .B1(_01774_),
    .B2(\i_exotiny._0018_[1] ),
    .A2(_01771_),
    .A1(\i_exotiny._0016_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05204_ (.Y(_01932_),
    .B1(_01783_),
    .B2(\i_exotiny._0023_[1] ),
    .A2(_01767_),
    .A1(\i_exotiny._0032_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05205_ (.B(_01926_),
    .C(_01931_),
    .A(_01924_),
    .Y(_01933_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01932_));
 sg13g2_nor2_1 _05206_ (.A(_01930_),
    .B(_01933_),
    .Y(_01934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05207_ (.Y(_01935_),
    .B1(_01791_),
    .B2(\i_exotiny._0026_[1] ),
    .A2(_01785_),
    .A1(\i_exotiny._0043_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05208_ (.Y(_01936_),
    .B1(_01790_),
    .B2(\i_exotiny._0034_[1] ),
    .A2(_01788_),
    .A1(\i_exotiny._0039_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05209_ (.B(_01921_),
    .C(_01935_),
    .A(_01755_),
    .Y(_01937_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01936_));
 sg13g2_a221oi_1 _05210_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0042_[1] ),
    .C1(_01937_),
    .B1(_01784_),
    .A1(\i_exotiny._0027_[1] ),
    .Y(_01938_),
    .A2(_01765_));
 sg13g2_a22oi_1 _05211_ (.Y(_01939_),
    .B1(_01772_),
    .B2(\i_exotiny._0033_[1] ),
    .A2(_01758_),
    .A1(\i_exotiny._0040_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05212_ (.B(_01927_),
    .C(_01939_),
    .A(_01922_),
    .Y(_01940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05213_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0038_[1] ),
    .C1(_01940_),
    .B1(_01792_),
    .A1(\i_exotiny._0014_[1] ),
    .Y(_01941_),
    .A2(_01760_));
 sg13g2_nand3_1 _05214_ (.B(_01938_),
    .C(_01941_),
    .A(_01934_),
    .Y(_01942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05215_ (.B1(_01942_),
    .VDD(VPWR),
    .Y(_01943_),
    .VSS(VGND),
    .A1(\i_exotiny._0036_[1] ),
    .A2(_01755_));
 sg13g2_a21oi_1 _05216_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01750_),
    .A2(_01943_),
    .Y(_01944_),
    .B1(net1108));
 sg13g2_a22oi_1 _05217_ (.Y(_01945_),
    .B1(_01920_),
    .B2(_01944_),
    .A2(net1108),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05218_ (.Y(_01946_),
    .B1(_01637_),
    .B2(\i_exotiny._0024_[1] ),
    .A2(_01636_),
    .A1(\i_exotiny._0019_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05219_ (.Y(_01947_),
    .B1(_01632_),
    .B2(\i_exotiny._0022_[1] ),
    .A2(_01628_),
    .A1(\i_exotiny._0037_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05220_ (.Y(_01948_),
    .B1(_01653_),
    .B2(\i_exotiny._0038_[1] ),
    .A2(_01618_),
    .A1(\i_exotiny._0031_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05221_ (.Y(_01949_),
    .B1(_01642_),
    .B2(\i_exotiny._0015_[1] ),
    .A2(_01638_),
    .A1(\i_exotiny._0029_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05222_ (.B(_01947_),
    .C(_01948_),
    .A(_01946_),
    .Y(_01950_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01949_));
 sg13g2_a22oi_1 _05223_ (.Y(_01951_),
    .B1(_01627_),
    .B2(\i_exotiny._0028_[1] ),
    .A2(_01622_),
    .A1(\i_exotiny._0023_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05224_ (.Y(_01952_),
    .B1(_01651_),
    .B2(\i_exotiny._0039_[1] ),
    .A2(_01621_),
    .A1(\i_exotiny._0043_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05225_ (.Y(_01953_),
    .B1(_01631_),
    .B2(\i_exotiny._0027_[1] ),
    .A2(_01626_),
    .A1(\i_exotiny._0014_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05226_ (.Y(_01954_),
    .B1(_01645_),
    .B2(\i_exotiny._0025_[1] ),
    .A2(_01625_),
    .A1(\i_exotiny._0030_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05227_ (.B(_01952_),
    .C(_01953_),
    .A(_01951_),
    .Y(_01955_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01954_));
 sg13g2_or2_1 _05228_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01956_),
    .B(\i_exotiny._0018_[1] ),
    .A(net1257));
 sg13g2_a22oi_1 _05229_ (.Y(_01957_),
    .B1(_01956_),
    .B2(_01643_),
    .A2(_01650_),
    .A1(\i_exotiny._0016_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05230_ (.Y(_01958_),
    .B1(_01649_),
    .B2(\i_exotiny._0042_[1] ),
    .A2(_01641_),
    .A1(\i_exotiny._0035_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05231_ (.Y(_01959_),
    .B1(_01648_),
    .B2(\i_exotiny._0033_[1] ),
    .A2(_01647_),
    .A1(\i_exotiny._0032_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05232_ (.Y(_01960_),
    .B1(_01624_),
    .B2(\i_exotiny._0040_[1] ),
    .A2(_01615_),
    .A1(\i_exotiny._0021_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05233_ (.Y(_01961_),
    .B1(_01630_),
    .B2(\i_exotiny._0041_[1] ),
    .A2(_01619_),
    .A1(\i_exotiny._0034_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05234_ (.Y(_01962_),
    .B1(_01655_),
    .B2(\i_exotiny._0026_[1] ),
    .A2(_01646_),
    .A1(\i_exotiny._0017_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05235_ (.Y(_01963_),
    .B1(_01654_),
    .B2(\i_exotiny._0020_[1] ),
    .A2(_01634_),
    .A1(\i_exotiny._0013_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _05236_ (.A(_01960_),
    .B(_01961_),
    .C(_01962_),
    .D(_01963_),
    .X(_01964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05237_ (.B(_01958_),
    .C(_01959_),
    .A(_01957_),
    .Y(_01965_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01964_));
 sg13g2_nor3_2 _05238_ (.A(_01950_),
    .B(_01955_),
    .C(_01965_),
    .Y(_01966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05239_ (.A(\i_exotiny._0036_[1] ),
    .B(_01644_),
    .Y(_01967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05240_ (.A(_01612_),
    .B(_01966_),
    .C(_01967_),
    .Y(_01968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05241_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ),
    .A2(_01612_),
    .Y(_01969_),
    .B1(_01968_));
 sg13g2_a221oi_1 _05242_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01944_),
    .C1(_01607_),
    .B1(_01920_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ),
    .Y(_01970_),
    .A2(net1107));
 sg13g2_and2_1 _05243_ (.A(net1110),
    .B(_01969_),
    .X(_01971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _05244_ (.A(_01970_),
    .B(_01971_),
    .Y(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05245_ (.A(_01825_),
    .B(_01970_),
    .C(_01971_),
    .Y(_01972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _05246_ (.Y(_01973_),
    .B(net35),
    .A_N(_01825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05247_ (.A(net1109),
    .B(_01969_),
    .X(_01974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05248_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01944_),
    .C1(net1109),
    .B1(_01920_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ),
    .Y(_01975_),
    .A2(net1107));
 sg13g2_nor2_1 _05249_ (.A(_01974_),
    .B(_01975_),
    .Y(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05250_ (.B1(_01831_),
    .VDD(VPWR),
    .Y(_01976_),
    .VSS(VGND),
    .A1(_01974_),
    .A2(_01975_));
 sg13g2_or3_1 _05251_ (.A(_01831_),
    .B(_01974_),
    .C(_01975_),
    .X(_01977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05252_ (.B(_01976_),
    .C(_01977_),
    .A(_01972_),
    .Y(_01978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _05253_ (.A2(_01977_),
    .A1(_01976_),
    .B1(_01972_),
    .X(_01979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05254_ (.Y(_01980_),
    .A(_01978_),
    .B(_01979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _05255_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01981_),
    .B(_01742_),
    .A(_01715_));
 sg13g2_a21oi_1 _05256_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01743_),
    .A2(_01981_),
    .Y(_01982_),
    .B1(_01702_));
 sg13g2_nand2_1 _05257_ (.Y(_01983_),
    .A(_01424_),
    .B(_01710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05258_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01371_),
    .A2(_01739_),
    .Y(_01984_),
    .B1(_01983_));
 sg13g2_a21o_1 _05259_ (.A2(_01983_),
    .A1(_01715_),
    .B1(_01701_),
    .X(_01985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05260_ (.B1(_01385_),
    .VDD(VPWR),
    .Y(_01986_),
    .VSS(VGND),
    .A1(_01984_),
    .A2(_01985_));
 sg13g2_a21oi_1 _05261_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1267),
    .A2(\i_exotiny._6090_[0] ),
    .Y(_01987_),
    .B1(_01750_));
 sg13g2_o21ai_1 _05262_ (.B1(_01987_),
    .VDD(VPWR),
    .Y(_01988_),
    .VSS(VGND),
    .A1(_01982_),
    .A2(_01986_));
 sg13g2_nand2_1 _05263_ (.Y(_01989_),
    .A(\i_exotiny._0015_[0] ),
    .B(_01761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05264_ (.Y(_01990_),
    .A(\i_exotiny._0023_[0] ),
    .B(_01783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05265_ (.Y(_01991_),
    .B1(_01777_),
    .B2(\i_exotiny._0013_[0] ),
    .A2(_01770_),
    .A1(\i_exotiny._0025_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05266_ (.Y(_01992_),
    .B1(_01781_),
    .B2(\i_exotiny._0028_[0] ),
    .A2(_01766_),
    .A1(\i_exotiny._0030_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05267_ (.Y(_01993_),
    .B1(_01787_),
    .B2(\i_exotiny._0031_[0] ),
    .A2(_01779_),
    .A1(\i_exotiny._0020_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05268_ (.Y(_01994_),
    .B1(_01786_),
    .B2(\i_exotiny._0017_[0] ),
    .A2(_01769_),
    .A1(\i_exotiny._0022_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05269_ (.Y(_01995_),
    .B1(_01776_),
    .B2(\i_exotiny._0021_[0] ),
    .A2(_01760_),
    .A1(\i_exotiny._0014_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05270_ (.B(_01993_),
    .C(_01994_),
    .A(_01991_),
    .Y(_01996_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01995_));
 sg13g2_a22oi_1 _05271_ (.Y(_01997_),
    .B1(_01792_),
    .B2(\i_exotiny._0038_[0] ),
    .A2(_01785_),
    .A1(\i_exotiny._0043_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05272_ (.Y(_01998_),
    .B1(_01791_),
    .B2(\i_exotiny._0026_[0] ),
    .A2(_01758_),
    .A1(\i_exotiny._0040_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05273_ (.B(_01992_),
    .C(_01997_),
    .A(_01990_),
    .Y(_01999_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01998_));
 sg13g2_nor2_1 _05274_ (.A(_01996_),
    .B(_01999_),
    .Y(_02000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05275_ (.Y(_02001_),
    .B1(_01789_),
    .B2(\i_exotiny._0024_[0] ),
    .A2(_01765_),
    .A1(\i_exotiny._0027_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05276_ (.Y(_02002_),
    .B1(_01790_),
    .B2(\i_exotiny._0034_[0] ),
    .A2(_01774_),
    .A1(\i_exotiny._0018_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05277_ (.B(_01989_),
    .C(_02001_),
    .A(_01755_),
    .Y(_02003_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02002_));
 sg13g2_a221oi_1 _05278_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0039_[0] ),
    .C1(_02003_),
    .B1(_01788_),
    .A1(\i_exotiny._0033_[0] ),
    .Y(_02004_),
    .A2(_01772_));
 sg13g2_a22oi_1 _05279_ (.Y(_02005_),
    .B1(_01780_),
    .B2(\i_exotiny._0041_[0] ),
    .A2(_01763_),
    .A1(\i_exotiny._0029_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05280_ (.Y(_02006_),
    .B1(_01784_),
    .B2(\i_exotiny._0042_[0] ),
    .A2(_01771_),
    .A1(\i_exotiny._0016_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05281_ (.Y(_02007_),
    .B1(_01778_),
    .B2(\i_exotiny._0035_[0] ),
    .A2(_01773_),
    .A1(\i_exotiny._0019_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05282_ (.B(_02006_),
    .C(_02007_),
    .A(_02005_),
    .Y(_02008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05283_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._0037_[0] ),
    .C1(_02008_),
    .B1(_01782_),
    .A1(\i_exotiny._0032_[0] ),
    .Y(_02009_),
    .A2(_01767_));
 sg13g2_nand3_1 _05284_ (.B(_02004_),
    .C(_02009_),
    .A(_02000_),
    .Y(_02010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05285_ (.B1(_02010_),
    .VDD(VPWR),
    .Y(_02011_),
    .VSS(VGND),
    .A1(\i_exotiny._0036_[0] ),
    .A2(_01755_));
 sg13g2_a21oi_1 _05286_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01750_),
    .A2(_02011_),
    .Y(_02012_),
    .B1(net1108));
 sg13g2_and2_1 _05287_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ),
    .B(net1107),
    .X(_02013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _05288_ (.A2(_02012_),
    .A1(_01988_),
    .B1(_02013_),
    .X(_02014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05289_ (.Y(_02015_),
    .B1(_01621_),
    .B2(\i_exotiny._0043_[0] ),
    .A2(_01619_),
    .A1(\i_exotiny._0034_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05290_ (.Y(_02016_),
    .B1(_01638_),
    .B2(\i_exotiny._0029_[0] ),
    .A2(_01626_),
    .A1(\i_exotiny._0014_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05291_ (.Y(_02017_),
    .B1(_01650_),
    .B2(\i_exotiny._0016_[0] ),
    .A2(_01641_),
    .A1(\i_exotiny._0035_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05292_ (.Y(_02018_),
    .B1(_01634_),
    .B2(\i_exotiny._0013_[0] ),
    .A2(_01627_),
    .A1(\i_exotiny._0028_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05293_ (.B(_02016_),
    .C(_02017_),
    .A(_02015_),
    .Y(_02019_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02018_));
 sg13g2_a22oi_1 _05294_ (.Y(_02020_),
    .B1(_01653_),
    .B2(\i_exotiny._0038_[0] ),
    .A2(_01642_),
    .A1(\i_exotiny._0015_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05295_ (.Y(_02021_),
    .B1(_01647_),
    .B2(\i_exotiny._0032_[0] ),
    .A2(_01645_),
    .A1(\i_exotiny._0025_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05296_ (.Y(_02022_),
    .B1(_01636_),
    .B2(\i_exotiny._0019_[0] ),
    .A2(_01628_),
    .A1(\i_exotiny._0037_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05297_ (.Y(_02023_),
    .B1(_01632_),
    .B2(\i_exotiny._0022_[0] ),
    .A2(_01622_),
    .A1(\i_exotiny._0023_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05298_ (.B(_02021_),
    .C(_02022_),
    .A(_02020_),
    .Y(_02024_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02023_));
 sg13g2_or2_1 _05299_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_02025_),
    .B(\i_exotiny._0018_[0] ),
    .A(net1257));
 sg13g2_a22oi_1 _05300_ (.Y(_02026_),
    .B1(_02025_),
    .B2(_01643_),
    .A2(_01646_),
    .A1(\i_exotiny._0017_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05301_ (.Y(_02027_),
    .B1(_01654_),
    .B2(\i_exotiny._0020_[0] ),
    .A2(_01618_),
    .A1(\i_exotiny._0031_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05302_ (.Y(_02028_),
    .B1(_01655_),
    .B2(\i_exotiny._0026_[0] ),
    .A2(_01651_),
    .A1(\i_exotiny._0039_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05303_ (.Y(_02029_),
    .B1(_01649_),
    .B2(\i_exotiny._0042_[0] ),
    .A2(_01625_),
    .A1(\i_exotiny._0030_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05304_ (.Y(_02030_),
    .B1(_01631_),
    .B2(\i_exotiny._0027_[0] ),
    .A2(_01624_),
    .A1(\i_exotiny._0040_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05305_ (.Y(_02031_),
    .B1(_01648_),
    .B2(\i_exotiny._0033_[0] ),
    .A2(_01637_),
    .A1(\i_exotiny._0024_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05306_ (.Y(_02032_),
    .B1(_01630_),
    .B2(\i_exotiny._0041_[0] ),
    .A2(_01615_),
    .A1(\i_exotiny._0021_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _05307_ (.A(_02029_),
    .B(_02030_),
    .C(_02031_),
    .D(_02032_),
    .X(_02033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05308_ (.B(_02027_),
    .C(_02028_),
    .A(_02026_),
    .Y(_02034_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02033_));
 sg13g2_nor3_2 _05309_ (.A(_02019_),
    .B(_02024_),
    .C(_02034_),
    .Y(_02035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05310_ (.A(\i_exotiny._0036_[0] ),
    .B(_01644_),
    .Y(_02036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05311_ (.A(_01612_),
    .B(_02035_),
    .C(_02036_),
    .Y(_02037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _05312_ (.A2(_01612_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ),
    .B1(_02037_),
    .X(_02038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05313_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02012_),
    .C1(net1110),
    .B1(_01988_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ),
    .Y(_02039_),
    .A2(net1107));
 sg13g2_nor2_1 _05314_ (.A(net1109),
    .B(_02038_),
    .Y(_02040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _05315_ (.A(_02039_),
    .B(_02040_),
    .Y(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _05316_ (.A(_01825_),
    .B(_02039_),
    .C(_02040_),
    .X(_02041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05317_ (.A(_01608_),
    .B(_02038_),
    .X(_02042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05318_ (.A(net1110),
    .B(_02038_),
    .Y(_02043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05319_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02012_),
    .C1(net1109),
    .B1(_01988_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ),
    .Y(_02044_),
    .A2(net1107));
 sg13g2_nor2_2 _05320_ (.A(_02043_),
    .B(_02044_),
    .Y(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05321_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net1110),
    .C1(_02042_),
    .B1(_02014_),
    .A1(\i_exotiny._0550_ ),
    .Y(_02045_),
    .A2(_01829_));
 sg13g2_nor3_1 _05322_ (.A(_01831_),
    .B(_02043_),
    .C(_02044_),
    .Y(_02046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05323_ (.A(_02045_),
    .B(_02046_),
    .Y(_02047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05324_ (.A(_02041_),
    .B(_02045_),
    .C(_02046_),
    .Y(_02048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _05325_ (.A(_02041_),
    .B(_02045_),
    .C(_02046_),
    .X(_02049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05326_ (.B1(_02041_),
    .VDD(VPWR),
    .Y(_02050_),
    .VSS(VGND),
    .A1(_02045_),
    .A2(_02046_));
 sg13g2_and2_1 _05327_ (.A(_02049_),
    .B(_02050_),
    .X(_02051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05328_ (.Y(_02052_),
    .B1(_02049_),
    .B2(_02050_),
    .A2(_01979_),
    .A1(_01978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05329_ (.A(\i_exotiny._0352_ ),
    .B(_01817_),
    .Y(_02053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05330_ (.B(_02052_),
    .C(_02053_),
    .A(_01912_),
    .Y(_02054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05331_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01388_),
    .A2(_02054_),
    .Y(_02055_),
    .B1(_01396_));
 sg13g2_o21ai_1 _05332_ (.B1(_01388_),
    .VDD(VPWR),
    .Y(_02056_),
    .VSS(VGND),
    .A1(\i_exotiny._0352_ ),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r ));
 sg13g2_nor2_1 _05333_ (.A(_01818_),
    .B(_02056_),
    .Y(_02057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _05334_ (.X(_02058_),
    .A(_01912_),
    .B(_02052_),
    .C(_02057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05335_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01976_),
    .A2(_01977_),
    .Y(_02059_),
    .B1(_01973_));
 sg13g2_a22oi_1 _05336_ (.Y(_02060_),
    .B1(_02041_),
    .B2(_02047_),
    .A2(_01979_),
    .A1(_01978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05337_ (.B1(_01912_),
    .VDD(VPWR),
    .Y(_02061_),
    .VSS(VGND),
    .A1(_02059_),
    .A2(_02060_));
 sg13g2_o21ai_1 _05338_ (.B1(\i_exotiny._1266_ ),
    .VDD(VPWR),
    .Y(_02062_),
    .VSS(VGND),
    .A1(_01459_),
    .A2(_01678_));
 sg13g2_nor2b_1 _05339_ (.A(_01828_),
    .B_N(_02062_),
    .Y(_02063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05340_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01832_),
    .A2(_01833_),
    .Y(_02064_),
    .B1(_02062_));
 sg13g2_or2_1 _05341_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_02065_),
    .B(_02064_),
    .A(_02063_));
 sg13g2_nand2_1 _05342_ (.Y(_02066_),
    .A(_01388_),
    .B(_01818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05343_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01905_),
    .A2(_01907_),
    .Y(_02067_),
    .B1(_01900_));
 sg13g2_a221oi_1 _05344_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01837_),
    .C1(_02066_),
    .B1(_02067_),
    .A1(_01834_),
    .Y(_02068_),
    .A2(_02065_));
 sg13g2_a21o_1 _05345_ (.A2(_02068_),
    .A1(_02061_),
    .B1(_02058_),
    .X(_02069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _05346_ (.VSS(VGND),
    .VDD(VPWR),
    .X(\i_exotiny._1207_ ),
    .B(_02069_),
    .A(_02055_));
 sg13g2_nand2b_1 _05347_ (.Y(_02070_),
    .B(net1116),
    .A_N(_01578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _05348_ (.B(\i_exotiny.i_wb_regs.spi_auto_cs_o ),
    .C(_02070_),
    .Y(_02071_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\i_exotiny.gpo[1] ));
 sg13g2_and2_1 _05349_ (.A(\i_exotiny.gpo[0] ),
    .B(_02071_),
    .X(gpo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05350_ (.A(net1263),
    .B(net3780),
    .Y(_02072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05351_ (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set [0]),
    .B_N(net1832),
    .Y(_02073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05352_ (.Y(_02074_),
    .A(net1263),
    .B(_01402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05353_ (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set [0]),
    .B(_02074_),
    .Y(_02075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _05354_ (.Y(_02076_),
    .B(net3326),
    .A_N(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05355_ (.Y(_02077_),
    .B1(_01400_),
    .B2(_01375_),
    .A2(\i_exotiny._2034_[1] ),
    .A1(_00015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _05356_ (.Y(_02078_),
    .A(_00018_),
    .B(\i_exotiny._2034_[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _05357_ (.B(\i_exotiny._2034_[8] ),
    .A(_00022_),
    .X(_02079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05358_ (.A(_00020_),
    .B(\i_exotiny._2034_[6] ),
    .Y(_02080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05359_ (.Y(_02081_),
    .A(_00020_),
    .B(\i_exotiny._2034_[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _05360_ (.B(\i_exotiny._2034_[9] ),
    .A(_00023_),
    .X(_02082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _05361_ (.B(\i_exotiny._2034_[5] ),
    .A(_00019_),
    .X(_02083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _05362_ (.B(\i_exotiny._2034_[3] ),
    .A(_00017_),
    .X(_02084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05363_ (.Y(_02085_),
    .B1(_01399_),
    .B2(_01376_),
    .A2(_01398_),
    .A1(_01377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05364_ (.Y(_02086_),
    .B1(\i_exotiny._2034_[7] ),
    .B2(_00021_),
    .A2(\i_exotiny._2034_[2] ),
    .A1(_00016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05365_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_00014_),
    .A2(\i_exotiny._2034_[0] ),
    .Y(_02087_),
    .B1(_02080_));
 sg13g2_nand4_1 _05366_ (.B(_02085_),
    .C(_02086_),
    .A(_02077_),
    .Y(_02088_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02087_));
 sg13g2_o21ai_1 _05367_ (.B1(_02081_),
    .VDD(VPWR),
    .Y(_02089_),
    .VSS(VGND),
    .A1(_00021_),
    .A2(\i_exotiny._2034_[7] ));
 sg13g2_nand4_1 _05368_ (.B(_02082_),
    .C(_02083_),
    .A(_02079_),
    .Y(_02090_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02084_));
 sg13g2_nor4_1 _05369_ (.A(_02078_),
    .B(_02088_),
    .C(_02089_),
    .D(_02090_),
    .Y(_02091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05370_ (.A(net1832),
    .B(_02076_),
    .C(net1112),
    .Y(_02092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05371_ (.A(net1263),
    .B(\i_exotiny.i_wdg_top.do_cnt ),
    .X(_02093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05372_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02092_),
    .A2(_02093_),
    .Y(_02094_),
    .B1(_02075_));
 sg13g2_nor2b_1 _05373_ (.A(net1832),
    .B_N(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.genblk7.g_value.r_value [0]),
    .Y(_02095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05374_ (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set [0]),
    .B(_02074_),
    .C(_02095_),
    .Y(_02096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05375_ (.A(net1263),
    .B(_01402_),
    .Y(_02097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05376_ (.A(net1263),
    .B(_01402_),
    .C(_02076_),
    .Y(_02098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05377_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1112),
    .A2(_02098_),
    .Y(_02099_),
    .B1(_02096_));
 sg13g2_nand2b_1 _05378_ (.Y(_02100_),
    .B(_02099_),
    .A_N(_02094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05379_ (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_hw_set [0]),
    .B(net3780),
    .C(_02076_),
    .Y(_02101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05380_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02092_),
    .A2(_02097_),
    .Y(_02102_),
    .B1(_02101_));
 sg13g2_a22oi_1 _05381_ (.Y(\i_exotiny._2055_[0] ),
    .B1(_02100_),
    .B2(_02102_),
    .A2(_02073_),
    .A1(net3781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _05382_ (.A2(_02093_),
    .A1(net1112),
    .B1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set [0]),
    .X(_02103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05383_ (.Y(_02104_),
    .A(_02073_),
    .B(_02093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05384_ (.B1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set [0]),
    .VDD(VPWR),
    .Y(_02105_),
    .VSS(VGND),
    .A1(net1832),
    .A2(_02074_));
 sg13g2_nand4_1 _05385_ (.B(_02103_),
    .C(_02104_),
    .A(net3326),
    .Y(_02106_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02105_));
 sg13g2_inv_1 _05386_ (.VDD(VPWR),
    .Y(\i_exotiny._2055_[2] ),
    .A(net3327),
    .VSS(VGND));
 sg13g2_a21oi_1 _05387_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02094_),
    .A2(_02106_),
    .Y(_02107_),
    .B1(_02096_));
 sg13g2_a21oi_1 _05388_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1112),
    .A2(_02098_),
    .Y(_02108_),
    .B1(_02107_));
 sg13g2_nor2_1 _05389_ (.A(net1832),
    .B(_02108_),
    .Y(\i_exotiny._2055_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05390_ (.A(\i_exotiny._2034_[0] ),
    .B(net1112),
    .Y(\i_exotiny._2043_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _05391_ (.Y(_02109_),
    .A(\i_exotiny._2034_[0] ),
    .B(\i_exotiny._2034_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05392_ (.A(net1112),
    .B(_02109_),
    .Y(\i_exotiny._2043_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05393_ (.B(\i_exotiny._2034_[1] ),
    .C(\i_exotiny._2034_[2] ),
    .A(\i_exotiny._2034_[0] ),
    .Y(_02110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05394_ (.B1(_01400_),
    .VDD(VPWR),
    .Y(_02111_),
    .VSS(VGND),
    .A1(_01398_),
    .A2(_01399_));
 sg13g2_nand2_1 _05395_ (.Y(_02112_),
    .A(_02110_),
    .B(_02111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05396_ (.A(net1112),
    .B(_02112_),
    .Y(\i_exotiny._2043_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05397_ (.A(_01401_),
    .B(_02110_),
    .Y(_02113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05398_ (.A(_01401_),
    .B(_02110_),
    .X(_02114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05399_ (.A(net1113),
    .B(_02113_),
    .C(_02114_),
    .Y(\i_exotiny._2043_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05400_ (.A(\i_exotiny._2034_[4] ),
    .B(_02113_),
    .X(_02115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05401_ (.A(\i_exotiny._2034_[4] ),
    .B(_02113_),
    .Y(_02116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05402_ (.A(net1113),
    .B(_02115_),
    .C(_02116_),
    .Y(\i_exotiny._2043_[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _05403_ (.Y(_02117_),
    .A(\i_exotiny._2034_[5] ),
    .B(_02115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05404_ (.A(net1112),
    .B(_02117_),
    .Y(\i_exotiny._2043_[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05405_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._2034_[5] ),
    .A2(_02115_),
    .Y(_02118_),
    .B1(\i_exotiny._2034_[6] ));
 sg13g2_and3_1 _05406_ (.X(_02119_),
    .A(\i_exotiny._2034_[5] ),
    .B(\i_exotiny._2034_[6] ),
    .C(_02115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05407_ (.A(net1113),
    .B(_02118_),
    .C(_02119_),
    .Y(\i_exotiny._2043_[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05408_ (.A(\i_exotiny._2034_[7] ),
    .B(_02119_),
    .Y(_02120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05409_ (.A(\i_exotiny._2034_[7] ),
    .B(_02119_),
    .X(_02121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05410_ (.A(net1113),
    .B(_02120_),
    .C(_02121_),
    .Y(\i_exotiny._2043_[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05411_ (.A(\i_exotiny._2034_[8] ),
    .B(_02121_),
    .Y(_02122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05412_ (.A(\i_exotiny._2034_[8] ),
    .B(_02121_),
    .X(_02123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05413_ (.A(net1113),
    .B(_02122_),
    .C(_02123_),
    .Y(\i_exotiny._2043_[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05414_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._2034_[9] ),
    .A2(_02123_),
    .Y(_02124_),
    .B1(net1113));
 sg13g2_o21ai_1 _05415_ (.B1(_02124_),
    .VDD(VPWR),
    .Y(_02125_),
    .VSS(VGND),
    .A1(\i_exotiny._2034_[9] ),
    .A2(_02123_));
 sg13g2_inv_1 _05416_ (.VDD(VPWR),
    .Y(\i_exotiny._2043_[9] ),
    .A(_02125_),
    .VSS(VGND));
 sg13g2_o21ai_1 _05417_ (.B1(_01529_),
    .VDD(VPWR),
    .Y(_02126_),
    .VSS(VGND),
    .A1(\i_exotiny._0327_[0] ),
    .A2(_01533_));
 sg13g2_nand3_1 _05418_ (.B(_01536_),
    .C(_02126_),
    .A(net1146),
    .Y(_02127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _05419_ (.B(_02127_),
    .A(\i_exotiny.i_wb_qspi_mem.cnt_r[2] ),
    .X(_02128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _05420_ (.VDD(VPWR),
    .Y(_02129_),
    .A(_02128_),
    .VSS(VGND));
 sg13g2_a21oi_1 _05421_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01387_),
    .A2(net1234),
    .Y(_02130_),
    .B1(net1244));
 sg13g2_nand3_1 _05422_ (.B(_01536_),
    .C(_02130_),
    .A(net1146),
    .Y(_02131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05423_ (.A(_01383_),
    .B(_02131_),
    .Y(_02132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _05424_ (.Y(_02133_),
    .A(net1230),
    .B(_02131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _05425_ (.Y(_02134_),
    .A(_01383_),
    .B(_02131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05426_ (.A(net1232),
    .B(_02129_),
    .C(_02134_),
    .Y(_02135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _05427_ (.A(_01384_),
    .B(_02134_),
    .Y(_02136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05428_ (.A(_01384_),
    .B(_02128_),
    .C(_02134_),
    .Y(_02137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _05429_ (.Y(_02138_),
    .A(_02129_),
    .B(_02136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05430_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1615_[0] ),
    .A2(_02136_),
    .Y(_02139_),
    .B1(_02137_));
 sg13g2_nor3_1 _05431_ (.A(net1232),
    .B(_02128_),
    .C(_02134_),
    .Y(_02140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05432_ (.Y(_02141_),
    .B1(_02140_),
    .B2(\i_exotiny._1618_[0] ),
    .A2(_02135_),
    .A1(\i_exotiny._1614_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _05433_ (.Y(_02142_),
    .A(_02128_),
    .B(_02132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _05434_ (.VDD(VPWR),
    .Y(_02143_),
    .A(_02142_),
    .VSS(VGND));
 sg13g2_nand2_1 _05435_ (.Y(_02144_),
    .A(net1232),
    .B(_02134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05436_ (.A(_02142_),
    .B(_02144_),
    .Y(_02145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05437_ (.A(net1232),
    .B(_02133_),
    .C(_02143_),
    .Y(_02146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05438_ (.Y(_02147_),
    .B1(_02146_),
    .B2(\i_exotiny._1616_[0] ),
    .A2(_02145_),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05439_ (.A(net1232),
    .B(_02133_),
    .C(_02142_),
    .Y(_02148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05440_ (.A(_02143_),
    .B(_02144_),
    .Y(_02149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05441_ (.Y(_02150_),
    .B1(_02149_),
    .B2(\i_exotiny._1617_[0] ),
    .A2(_02148_),
    .A1(\i_exotiny._1612_[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05442_ (.B(_02141_),
    .C(_02147_),
    .A(_02139_),
    .Y(_02151_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02150_));
 sg13g2_o21ai_1 _05443_ (.B1(net1264),
    .VDD(VPWR),
    .Y(_02152_),
    .VSS(VGND),
    .A1(\i_exotiny._1619_[0] ),
    .A2(_02138_));
 sg13g2_nand2b_1 _05444_ (.Y(_02153_),
    .B(_02151_),
    .A_N(_02152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05445_ (.B1(_02153_),
    .VDD(VPWR),
    .Y(net27),
    .VSS(VGND),
    .A1(\i_exotiny._1660_ ),
    .A2(_01403_));
 sg13g2_nand2b_1 _05446_ (.Y(_02154_),
    .B(\i_exotiny._0369_[5] ),
    .A_N(net1264),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05447_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1615_[1] ),
    .A2(_02136_),
    .Y(_02155_),
    .B1(_02137_));
 sg13g2_a22oi_1 _05448_ (.Y(_02156_),
    .B1(_02140_),
    .B2(\i_exotiny._1618_[1] ),
    .A2(_02135_),
    .A1(\i_exotiny._1614_[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05449_ (.Y(_02157_),
    .B1(_02146_),
    .B2(\i_exotiny._1616_[1] ),
    .A2(_02145_),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05450_ (.B(_02156_),
    .C(_02157_),
    .A(_02155_),
    .Y(_02158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05451_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._1617_[1] ),
    .C1(_02158_),
    .B1(_02149_),
    .A1(\i_exotiny._1612_[1] ),
    .Y(_02159_),
    .A2(_02148_));
 sg13g2_o21ai_1 _05452_ (.B1(net1264),
    .VDD(VPWR),
    .Y(_02160_),
    .VSS(VGND),
    .A1(\i_exotiny._1619_[1] ),
    .A2(_02138_));
 sg13g2_o21ai_1 _05453_ (.B1(_02154_),
    .VDD(VPWR),
    .Y(net28),
    .VSS(VGND),
    .A1(_02159_),
    .A2(_02160_));
 sg13g2_a21o_1 _05454_ (.A2(_02136_),
    .A1(\i_exotiny._1615_[2] ),
    .B1(_02137_),
    .X(_02161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05455_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._1618_[2] ),
    .C1(_02161_),
    .B1(_02140_),
    .A1(\i_exotiny._1614_[2] ),
    .Y(_02162_),
    .A2(_02135_));
 sg13g2_a22oi_1 _05456_ (.Y(_02163_),
    .B1(_02146_),
    .B2(\i_exotiny._1616_[2] ),
    .A2(_02145_),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05457_ (.Y(_02164_),
    .B1(_02149_),
    .B2(\i_exotiny._1617_[2] ),
    .A2(_02148_),
    .A1(\i_exotiny._1612_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05458_ (.B(_02163_),
    .C(_02164_),
    .A(_02162_),
    .Y(_02165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05459_ (.B1(\i_exotiny._1660_ ),
    .VDD(VPWR),
    .Y(_02166_),
    .VSS(VGND),
    .A1(\i_exotiny._1619_[2] ),
    .A2(_02138_));
 sg13g2_nand2b_1 _05460_ (.Y(_02167_),
    .B(_02165_),
    .A_N(_02166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05461_ (.B1(_02167_),
    .VDD(VPWR),
    .Y(net30),
    .VSS(VGND),
    .A1(net1264),
    .A2(_01404_));
 sg13g2_nand2b_1 _05462_ (.Y(_02168_),
    .B(\i_exotiny._0369_[7] ),
    .A_N(net1264),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05463_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1615_[3] ),
    .A2(_02136_),
    .Y(_02169_),
    .B1(_02137_));
 sg13g2_a22oi_1 _05464_ (.Y(_02170_),
    .B1(_02140_),
    .B2(\i_exotiny._1618_[3] ),
    .A2(_02135_),
    .A1(\i_exotiny._1614_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05465_ (.Y(_02171_),
    .B1(_02149_),
    .B2(\i_exotiny._1617_[3] ),
    .A2(_02148_),
    .A1(\i_exotiny._1612_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05466_ (.B(_02170_),
    .C(_02171_),
    .A(_02169_),
    .Y(_02172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05467_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\i_exotiny._1616_[3] ),
    .C1(_02172_),
    .B1(_02146_),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data [0]),
    .Y(_02173_),
    .A2(_02145_));
 sg13g2_o21ai_1 _05468_ (.B1(net1264),
    .VDD(VPWR),
    .Y(_02174_),
    .VSS(VGND),
    .A1(\i_exotiny._1619_[3] ),
    .A2(_02138_));
 sg13g2_o21ai_1 _05469_ (.B1(_02168_),
    .VDD(VPWR),
    .Y(net31),
    .VSS(VGND),
    .A1(_02173_),
    .A2(_02174_));
 sg13g2_and3_1 _05470_ (.X(\i_exotiny._1611_[1] ),
    .A(net1281),
    .B(net3702),
    .C(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05471_ (.B1(net1076),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[2] ),
    .VSS(VGND),
    .A1(_01405_),
    .A2(_01543_));
 sg13g2_and3_1 _05472_ (.X(\i_exotiny._1611_[3] ),
    .A(net1281),
    .B(net3702),
    .C(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05473_ (.A(net1265),
    .B(\i_exotiny._1711_ ),
    .C(_01521_),
    .Y(_02175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05474_ (.Y(_02176_),
    .A(net1284),
    .B(net3594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05475_ (.B1(net1076),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[5] ),
    .VSS(VGND),
    .A1(_02175_),
    .A2(_02176_));
 sg13g2_a21o_1 _05476_ (.A2(_01511_),
    .A1(net1265),
    .B1(_01545_),
    .X(_02177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _05477_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_02178_),
    .B(\i_exotiny._1757_ ),
    .A(net1265));
 sg13g2_nor2_1 _05478_ (.A(net3707),
    .B(_02177_),
    .Y(_02179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05479_ (.Y(_02180_),
    .A(_02178_),
    .B(_02179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _05480_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net1225),
    .Y(_02181_),
    .A2(_02179_),
    .A1(_02178_));
 sg13g2_and2_1 _05481_ (.A(net1872),
    .B(net1070),
    .X(\i_exotiny._1611_[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05482_ (.Y(_02182_),
    .A(net1284),
    .B(net3584),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05483_ (.B1(net1076),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[7] ),
    .VSS(VGND),
    .A1(_02175_),
    .A2(_02182_));
 sg13g2_nand2_1 _05484_ (.Y(_02183_),
    .A(net1283),
    .B(_01512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05485_ (.Y(_02184_),
    .A(net3601),
    .B(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05486_ (.B1(_02184_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[9] ),
    .VSS(VGND),
    .A1(_02127_),
    .A2(_02183_));
 sg13g2_nand2_1 _05487_ (.Y(_02185_),
    .A(net3457),
    .B(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05488_ (.A(net1279),
    .B_N(net1233),
    .Y(_02186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05489_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0314_[2] ),
    .A2(net1277),
    .Y(_02187_),
    .B1(_02186_));
 sg13g2_o21ai_1 _05490_ (.B1(_02185_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[10] ),
    .VSS(VGND),
    .A1(net1074),
    .A2(_02187_));
 sg13g2_nand2_1 _05491_ (.Y(_02188_),
    .A(net3387),
    .B(net1070),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05492_ (.A(net1274),
    .B(_01390_),
    .Y(_02189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05493_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0314_[3] ),
    .A2(net1279),
    .Y(_02190_),
    .B1(_02189_));
 sg13g2_o21ai_1 _05494_ (.B1(_02188_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[11] ),
    .VSS(VGND),
    .A1(net1075),
    .A2(_02190_));
 sg13g2_nand2_1 _05495_ (.Y(_02191_),
    .A(net3675),
    .B(net1070),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05496_ (.A(net1279),
    .B(_01393_),
    .Y(_02192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05497_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3603),
    .A2(net1279),
    .Y(_02193_),
    .B1(_02192_));
 sg13g2_o21ai_1 _05498_ (.B1(_02191_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[13] ),
    .VSS(VGND),
    .A1(net1076),
    .A2(_02193_));
 sg13g2_nand2_1 _05499_ (.Y(_02194_),
    .A(net3737),
    .B(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05500_ (.A(net1278),
    .B(_01386_),
    .Y(_02195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05501_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3407),
    .A2(net1276),
    .Y(_02196_),
    .B1(_02195_));
 sg13g2_o21ai_1 _05502_ (.B1(_02194_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[14] ),
    .VSS(VGND),
    .A1(net1074),
    .A2(_02196_));
 sg13g2_nand2_1 _05503_ (.Y(_02197_),
    .A(net3505),
    .B(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05504_ (.A(net1280),
    .B_N(\i_exotiny._0315_[7] ),
    .Y(_02198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05505_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0314_[7] ),
    .A2(net1280),
    .Y(_02199_),
    .B1(_02198_));
 sg13g2_o21ai_1 _05506_ (.B1(_02197_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[15] ),
    .VSS(VGND),
    .A1(net1074),
    .A2(_02199_));
 sg13g2_nand2_1 _05507_ (.Y(_02200_),
    .A(net2125),
    .B(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05508_ (.A(net1275),
    .B_N(\i_exotiny._0315_[9] ),
    .Y(_02201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05509_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0314_[9] ),
    .A2(net1275),
    .Y(_02202_),
    .B1(_02201_));
 sg13g2_o21ai_1 _05510_ (.B1(_02200_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[17] ),
    .VSS(VGND),
    .A1(net1074),
    .A2(_02202_));
 sg13g2_nand2_1 _05511_ (.Y(_02203_),
    .A(net3307),
    .B(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05512_ (.A(net1276),
    .B_N(\i_exotiny._0315_[10] ),
    .Y(_02204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05513_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0314_[10] ),
    .A2(net1276),
    .Y(_02205_),
    .B1(_02204_));
 sg13g2_o21ai_1 _05514_ (.B1(_02203_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[18] ),
    .VSS(VGND),
    .A1(net1074),
    .A2(_02205_));
 sg13g2_nand2_1 _05515_ (.Y(_02206_),
    .A(net2061),
    .B(net1070),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05516_ (.A(net1277),
    .B_N(\i_exotiny._0315_[11] ),
    .Y(_02207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05517_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0314_[11] ),
    .A2(net1276),
    .Y(_02208_),
    .B1(_02207_));
 sg13g2_o21ai_1 _05518_ (.B1(_02206_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[19] ),
    .VSS(VGND),
    .A1(net1075),
    .A2(_02208_));
 sg13g2_nand2_1 _05519_ (.Y(_02209_),
    .A(net2997),
    .B(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05520_ (.A(net1275),
    .B_N(\i_exotiny._0315_[13] ),
    .Y(_02210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05521_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0314_[13] ),
    .A2(net1275),
    .Y(_02211_),
    .B1(_02210_));
 sg13g2_o21ai_1 _05522_ (.B1(_02209_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[21] ),
    .VSS(VGND),
    .A1(net1074),
    .A2(_02211_));
 sg13g2_nand2_1 _05523_ (.Y(_02212_),
    .A(net3443),
    .B(net1070),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05524_ (.A(net1276),
    .B_N(\i_exotiny._0315_[14] ),
    .Y(_02213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05525_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0314_[14] ),
    .A2(net1276),
    .Y(_02214_),
    .B1(_02213_));
 sg13g2_o21ai_1 _05526_ (.B1(_02212_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[22] ),
    .VSS(VGND),
    .A1(net1075),
    .A2(_02214_));
 sg13g2_nand2_1 _05527_ (.Y(_02215_),
    .A(net3641),
    .B(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05528_ (.A(net1277),
    .B_N(net3612),
    .Y(_02216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05529_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3498),
    .A2(net1276),
    .Y(_02217_),
    .B1(_02216_));
 sg13g2_o21ai_1 _05530_ (.B1(_02215_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[23] ),
    .VSS(VGND),
    .A1(net1075),
    .A2(_02217_));
 sg13g2_nand2_1 _05531_ (.Y(_02218_),
    .A(net3749),
    .B(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05532_ (.B1(net1284),
    .VDD(VPWR),
    .Y(_02219_),
    .VSS(VGND),
    .A1(\i_exotiny._1711_ ),
    .A2(_02178_));
 sg13g2_and2_1 _05533_ (.A(net1218),
    .B(_01520_),
    .X(_02220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05534_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_wb_qspi_mem.crm_r ),
    .A2(_01520_),
    .Y(_02221_),
    .B1(_01512_));
 sg13g2_nand2_1 _05535_ (.Y(_02222_),
    .A(net2864),
    .B(net1272),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _05536_ (.Y(_02223_),
    .B(net3706),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1272));
 sg13g2_a221oi_1 _05537_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02223_),
    .C1(_02221_),
    .B1(_02222_),
    .A1(_01484_),
    .Y(_02224_),
    .A2(_01513_));
 sg13g2_a21oi_1 _05538_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01485_),
    .A2(_02220_),
    .Y(_02225_),
    .B1(_02224_));
 sg13g2_nor2_1 _05539_ (.A(\i_exotiny.i_wb_qspi_mem.crm_r ),
    .B(net1218),
    .Y(_02226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05540_ (.B1(_02218_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[25] ),
    .VSS(VGND),
    .A1(_02219_),
    .A2(_02225_));
 sg13g2_nand2_1 _05541_ (.Y(_02227_),
    .A(net3643),
    .B(net1070),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05542_ (.A(net1277),
    .B_N(net3549),
    .Y(_02228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05543_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3402),
    .A2(net1276),
    .Y(_02229_),
    .B1(_02228_));
 sg13g2_o21ai_1 _05544_ (.B1(_02227_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[26] ),
    .VSS(VGND),
    .A1(net1074),
    .A2(_02229_));
 sg13g2_nand2_1 _05545_ (.Y(_02230_),
    .A(net3596),
    .B(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _05546_ (.Y(_02231_),
    .B(net1275),
    .A_N(\i_exotiny._0314_[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05547_ (.B1(_02231_),
    .VDD(VPWR),
    .Y(_02232_),
    .VSS(VGND),
    .A1(net1275),
    .A2(\i_exotiny._0315_[19] ));
 sg13g2_nor2_1 _05548_ (.A(_02221_),
    .B(_02232_),
    .Y(_02233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05549_ (.A(_01553_),
    .B(_02220_),
    .C(_02233_),
    .Y(_02234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05550_ (.B1(_02230_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[27] ),
    .VSS(VGND),
    .A1(_02219_),
    .A2(_02234_));
 sg13g2_nand2_1 _05551_ (.Y(_02235_),
    .A(net2735),
    .B(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05552_ (.A0(\i_exotiny._0315_[21] ),
    .A1(\i_exotiny._0314_[21] ),
    .S(net1272),
    .X(_02236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05553_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01523_),
    .A2(_02236_),
    .Y(_02237_),
    .B1(_01553_));
 sg13g2_o21ai_1 _05554_ (.B1(_02235_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[29] ),
    .VSS(VGND),
    .A1(_02219_),
    .A2(_02237_));
 sg13g2_nand2_1 _05555_ (.Y(_02238_),
    .A(net3798),
    .B(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05556_ (.A(net1277),
    .B_N(\i_exotiny._0315_[22] ),
    .Y(_02239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05557_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3610),
    .A2(net1277),
    .Y(_02240_),
    .B1(_02239_));
 sg13g2_o21ai_1 _05558_ (.B1(_02238_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[30] ),
    .VSS(VGND),
    .A1(net1074),
    .A2(_02240_));
 sg13g2_nand2_1 _05559_ (.Y(_02241_),
    .A(net3729),
    .B(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05560_ (.A(net1275),
    .B_N(net3185),
    .Y(_02242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05561_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3155),
    .A2(net1275),
    .Y(_02243_),
    .B1(_02242_));
 sg13g2_o21ai_1 _05562_ (.B1(_02241_),
    .VDD(VPWR),
    .Y(\i_exotiny._1611_[31] ),
    .VSS(VGND),
    .A1(net1076),
    .A2(_02243_));
 sg13g2_xnor2_1 _05563_ (.Y(_02244_),
    .A(\i_exotiny._0315_[7] ),
    .B(_01690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05564_ (.A(\i_exotiny._0327_[0] ),
    .B(net1201),
    .Y(_02245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05565_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1202),
    .A2(_02244_),
    .Y(_02246_),
    .B1(_02245_));
 sg13g2_o21ai_1 _05566_ (.B1(net1266),
    .VDD(VPWR),
    .Y(_02247_),
    .VSS(VGND),
    .A1(net3523),
    .A2(net3677));
 sg13g2_a21oi_1 _05567_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3523),
    .A2(net3677),
    .Y(_02248_),
    .B1(_02247_));
 sg13g2_a21oi_1 _05568_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01385_),
    .A2(_02246_),
    .Y(\i_exotiny._1489_[1] ),
    .B1(net3678));
 sg13g2_o21ai_1 _05569_ (.B1(_01424_),
    .VDD(VPWR),
    .Y(_02249_),
    .VSS(VGND),
    .A1(\i_exotiny._0315_[7] ),
    .A2(\i_exotiny._0315_[6] ));
 sg13g2_xnor2_1 _05570_ (.Y(_02250_),
    .A(\i_exotiny._0315_[8] ),
    .B(_02249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _05571_ (.B(net1234),
    .A(\i_exotiny._0327_[0] ),
    .X(_02251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05572_ (.A(net1201),
    .B(_02251_),
    .Y(_02252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05573_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1202),
    .A2(_02250_),
    .Y(_02253_),
    .B1(_02252_));
 sg13g2_o21ai_1 _05574_ (.B1(net1984),
    .VDD(VPWR),
    .Y(_02254_),
    .VSS(VGND),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0] ),
    .A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1] ));
 sg13g2_nor2_1 _05575_ (.A(_01385_),
    .B(_01439_),
    .Y(_02255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05576_ (.Y(\i_exotiny._1489_[2] ),
    .B1(net1985),
    .B2(_02255_),
    .A2(_02253_),
    .A1(_01385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05577_ (.Y(_02256_),
    .A(net2570),
    .B(net1291),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _05578_ (.A(net1204),
    .Y(\i_exotiny._0000_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05579_ (.A(net1197),
    .B(net1212),
    .Y(_00000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _05580_ (.A(\i_exotiny._1793_ ),
    .B(net1218),
    .C(_01555_),
    .X(\i_exotiny._5420_$func$/home/user/heichips25-fazyrv-exotiny/build/exotiny_preproc.v:7404$13.$result [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05581_ (.A(_01402_),
    .B(net1204),
    .Y(\i_exotiny._2032_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _05582_ (.B(_01465_),
    .C(net1201),
    .Y(_02257_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_01461_));
 sg13g2_nand3_1 _05583_ (.B(\i_exotiny._0352_ ),
    .C(_02257_),
    .A(net1269),
    .Y(_02258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05584_ (.B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ),
    .C(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r [0]),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ),
    .Y(_02259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05585_ (.Y(_02260_),
    .A(\i_exotiny._1306_ ),
    .B(\i_exotiny._0352_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05586_ (.B1(_02259_),
    .VDD(VPWR),
    .Y(_02261_),
    .VSS(VGND),
    .A1(_02257_),
    .A2(_02260_));
 sg13g2_nor2b_1 _05587_ (.A(_02261_),
    .B_N(_02258_),
    .Y(_02262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05588_ (.A(_02262_),
    .B_N(\i_exotiny._0314_[2] ),
    .Y(_02263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05589_ (.A(net3390),
    .B(_02263_),
    .X(\i_exotiny._1465_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05590_ (.A(\i_exotiny._0352_ ),
    .B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r ),
    .Y(_02264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05591_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0352_ ),
    .A2(_01831_),
    .Y(_02265_),
    .B1(_02264_));
 sg13g2_a21oi_1 _05592_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02050_),
    .A2(_02265_),
    .Y(_02266_),
    .B1(_02048_));
 sg13g2_o21ai_1 _05593_ (.B1(_01978_),
    .VDD(VPWR),
    .Y(_02267_),
    .VSS(VGND),
    .A1(_01980_),
    .A2(_02266_));
 sg13g2_a21oi_1 _05594_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01911_),
    .A2(_02267_),
    .Y(_02268_),
    .B1(_01909_));
 sg13g2_a21o_1 _05595_ (.A2(_02267_),
    .A1(_01911_),
    .B1(_01909_),
    .X(_02269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05596_ (.B1(_01834_),
    .VDD(VPWR),
    .Y(\i_exotiny._1206_ ),
    .VSS(VGND),
    .A1(_01837_),
    .A2(_02268_));
 sg13g2_nor2_1 _05597_ (.A(_01473_),
    .B(_02260_),
    .Y(ccx_req),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05598_ (.A(net3326),
    .B(net1105),
    .Y(_02270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05599_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01361_),
    .A2(net1105),
    .Y(_00024_),
    .B1(_02270_));
 sg13g2_nor2_1 _05600_ (.A(net3511),
    .B(net1105),
    .Y(_02271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05601_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1612_[0] ),
    .A2(net1106),
    .Y(_00025_),
    .B1(_02271_));
 sg13g2_nor2_1 _05602_ (.A(\i_exotiny._1956_ ),
    .B(_01571_),
    .Y(_02272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05603_ (.A(net1072),
    .B(_02272_),
    .Y(_02273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05604_ (.A(net1978),
    .B(net1060),
    .Y(_02274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05605_ (.A0(_01397_),
    .A1(_01366_),
    .S(net1116),
    .X(_02275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05606_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1060),
    .A2(_02275_),
    .Y(_00027_),
    .B1(_02274_));
 sg13g2_nor2b_1 _05607_ (.A(net1116),
    .B_N(\i_exotiny._1924_[2] ),
    .Y(_02276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05608_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data [0]),
    .A2(net1118),
    .Y(_02277_),
    .B1(_02276_));
 sg13g2_nor2_1 _05609_ (.A(net1903),
    .B(net1067),
    .Y(_02278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05610_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1067),
    .A2(_02277_),
    .Y(_00028_),
    .B1(_02278_));
 sg13g2_nor2_1 _05611_ (.A(net1907),
    .B(net1061),
    .Y(_02279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05612_ (.A(net1119),
    .B_N(net1903),
    .Y(_02280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05613_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data [0]),
    .A2(net1119),
    .Y(_02281_),
    .B1(_02280_));
 sg13g2_a21oi_1 _05614_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1067),
    .A2(_02281_),
    .Y(_00029_),
    .B1(_02279_));
 sg13g2_nor2_1 _05615_ (.A(net2050),
    .B(net1061),
    .Y(_02282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05616_ (.A(net1120),
    .B_N(net1907),
    .Y(_02283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05617_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1612_[0] ),
    .A2(net1119),
    .Y(_02284_),
    .B1(_02283_));
 sg13g2_a21oi_1 _05618_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1061),
    .A2(_02284_),
    .Y(_00030_),
    .B1(_02282_));
 sg13g2_nor2_1 _05619_ (.A(net1987),
    .B(net1065),
    .Y(_02285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05620_ (.A(net1119),
    .B_N(\i_exotiny._1924_[5] ),
    .Y(_02286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05621_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1612_[1] ),
    .A2(net1120),
    .Y(_02287_),
    .B1(_02286_));
 sg13g2_a21oi_1 _05622_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1061),
    .A2(_02287_),
    .Y(_00031_),
    .B1(_02285_));
 sg13g2_nor2_1 _05623_ (.A(net1895),
    .B(net1065),
    .Y(_02288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05624_ (.A(net1125),
    .B_N(\i_exotiny._1924_[6] ),
    .Y(_02289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05625_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1612_[2] ),
    .A2(net1124),
    .Y(_02290_),
    .B1(_02289_));
 sg13g2_a21oi_1 _05626_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1066),
    .A2(_02290_),
    .Y(_00032_),
    .B1(_02288_));
 sg13g2_nor2b_1 _05627_ (.A(net1124),
    .B_N(net1895),
    .Y(_02291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05628_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1612_[3] ),
    .A2(net1124),
    .Y(_02292_),
    .B1(_02291_));
 sg13g2_nor2_1 _05629_ (.A(net1941),
    .B(net1065),
    .Y(_02293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1065),
    .A2(_02292_),
    .Y(_00033_),
    .B1(_02293_));
 sg13g2_nor2_1 _05631_ (.A(net1943),
    .B(net1065),
    .Y(_02294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05632_ (.A(net1124),
    .B_N(net1941),
    .Y(_02295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05633_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1615_[0] ),
    .A2(net1125),
    .Y(_02296_),
    .B1(_02295_));
 sg13g2_a21oi_1 _05634_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1066),
    .A2(_02296_),
    .Y(_00034_),
    .B1(_02294_));
 sg13g2_nor2_1 _05635_ (.A(net2006),
    .B(net1065),
    .Y(_02297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05636_ (.A(net1119),
    .B_N(net1943),
    .Y(_02298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05637_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1615_[1] ),
    .A2(net1119),
    .Y(_02299_),
    .B1(_02298_));
 sg13g2_a21oi_1 _05638_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1061),
    .A2(_02299_),
    .Y(_00035_),
    .B1(_02297_));
 sg13g2_nor2_1 _05639_ (.A(net1909),
    .B(net1065),
    .Y(_02300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05640_ (.A(net1124),
    .B_N(\i_exotiny._1924_[10] ),
    .Y(_02301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05641_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1615_[2] ),
    .A2(net1124),
    .Y(_02302_),
    .B1(_02301_));
 sg13g2_a21oi_1 _05642_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1065),
    .A2(_02302_),
    .Y(_00036_),
    .B1(_02300_));
 sg13g2_nor2_1 _05643_ (.A(net1922),
    .B(net1066),
    .Y(_02303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05644_ (.A(net1124),
    .B_N(net1909),
    .Y(_02304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05645_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1615_[3] ),
    .A2(net1124),
    .Y(_02305_),
    .B1(_02304_));
 sg13g2_a21oi_1 _05646_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1066),
    .A2(_02305_),
    .Y(_00037_),
    .B1(_02303_));
 sg13g2_nor2b_1 _05647_ (.A(net1125),
    .B_N(net1922),
    .Y(_02306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05648_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1614_[0] ),
    .A2(net1125),
    .Y(_02307_),
    .B1(_02306_));
 sg13g2_nor2_1 _05649_ (.A(net1953),
    .B(net1066),
    .Y(_02308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05650_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1066),
    .A2(_02307_),
    .Y(_00038_),
    .B1(_02308_));
 sg13g2_nor2_1 _05651_ (.A(net1939),
    .B(net1066),
    .Y(_02309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05652_ (.A(net1125),
    .B_N(\i_exotiny._1924_[13] ),
    .Y(_02310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05653_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1614_[1] ),
    .A2(net1125),
    .Y(_02311_),
    .B1(_02310_));
 sg13g2_a21oi_1 _05654_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1067),
    .A2(_02311_),
    .Y(_00039_),
    .B1(_02309_));
 sg13g2_nor2_1 _05655_ (.A(net1963),
    .B(net1063),
    .Y(_02312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05656_ (.A(net1122),
    .B_N(net1939),
    .Y(_02313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05657_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1614_[2] ),
    .A2(net1122),
    .Y(_02314_),
    .B1(_02313_));
 sg13g2_a21oi_1 _05658_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1063),
    .A2(_02314_),
    .Y(_00040_),
    .B1(_02312_));
 sg13g2_nor2_1 _05659_ (.A(net2004),
    .B(net1063),
    .Y(_02315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05660_ (.A(net1122),
    .B_N(net1963),
    .Y(_02316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05661_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1614_[3] ),
    .A2(net1122),
    .Y(_02317_),
    .B1(_02316_));
 sg13g2_a21oi_1 _05662_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1063),
    .A2(_02317_),
    .Y(_00041_),
    .B1(_02315_));
 sg13g2_nor2b_1 _05663_ (.A(net1122),
    .B_N(net2004),
    .Y(_02318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05664_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1617_[0] ),
    .A2(net1123),
    .Y(_02319_),
    .B1(_02318_));
 sg13g2_nor2_1 _05665_ (.A(net2031),
    .B(net1064),
    .Y(_02320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05666_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1064),
    .A2(_02319_),
    .Y(_00042_),
    .B1(_02320_));
 sg13g2_nor2_1 _05667_ (.A(net1901),
    .B(net1062),
    .Y(_02321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05668_ (.A(net1123),
    .B_N(\i_exotiny._1924_[17] ),
    .Y(_02322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05669_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1617_[1] ),
    .A2(net1122),
    .Y(_02323_),
    .B1(_02322_));
 sg13g2_a21oi_1 _05670_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1062),
    .A2(_02323_),
    .Y(_00043_),
    .B1(_02321_));
 sg13g2_nor2_1 _05671_ (.A(net1947),
    .B(net1062),
    .Y(_02324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05672_ (.A(net1123),
    .B_N(net1901),
    .Y(_02325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05673_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1617_[2] ),
    .A2(net1121),
    .Y(_02326_),
    .B1(_02325_));
 sg13g2_a21oi_1 _05674_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1062),
    .A2(_02326_),
    .Y(_00044_),
    .B1(_02324_));
 sg13g2_nor2_1 _05675_ (.A(net1957),
    .B(net1062),
    .Y(_02327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05676_ (.A(net1121),
    .B_N(net1947),
    .Y(_02328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05677_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1617_[3] ),
    .A2(net1121),
    .Y(_02329_),
    .B1(_02328_));
 sg13g2_a21oi_1 _05678_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1062),
    .A2(_02329_),
    .Y(_00045_),
    .B1(_02327_));
 sg13g2_nor2_1 _05679_ (.A(net1916),
    .B(net1062),
    .Y(_02330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05680_ (.A(net1121),
    .B_N(\i_exotiny._1924_[20] ),
    .Y(_02331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05681_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1616_[0] ),
    .A2(net1121),
    .Y(_02332_),
    .B1(_02331_));
 sg13g2_a21oi_1 _05682_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1063),
    .A2(_02332_),
    .Y(_00046_),
    .B1(_02330_));
 sg13g2_nor2_1 _05683_ (.A(net1926),
    .B(net1063),
    .Y(_02333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05684_ (.A(net1121),
    .B_N(net1916),
    .Y(_02334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05685_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1616_[1] ),
    .A2(net1121),
    .Y(_02335_),
    .B1(_02334_));
 sg13g2_a21oi_1 _05686_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1063),
    .A2(_02335_),
    .Y(_00047_),
    .B1(_02333_));
 sg13g2_nor2_1 _05687_ (.A(net2046),
    .B(net1064),
    .Y(_02336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05688_ (.A(net1122),
    .B_N(net1926),
    .Y(_02337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05689_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1616_[2] ),
    .A2(net1121),
    .Y(_02338_),
    .B1(_02337_));
 sg13g2_a21oi_1 _05690_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1062),
    .A2(_02338_),
    .Y(_00048_),
    .B1(_02336_));
 sg13g2_nor2b_1 _05691_ (.A(net1123),
    .B_N(net2046),
    .Y(_02339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05692_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1616_[3] ),
    .A2(net1123),
    .Y(_02340_),
    .B1(_02339_));
 sg13g2_nor2_1 _05693_ (.A(net2528),
    .B(net1064),
    .Y(_02341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05694_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1064),
    .A2(_02340_),
    .Y(_00049_),
    .B1(_02341_));
 sg13g2_nor2_1 _05695_ (.A(net1920),
    .B(net1061),
    .Y(_02342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05696_ (.A(net1117),
    .B_N(\i_exotiny._1924_[24] ),
    .Y(_02343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05697_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1619_[0] ),
    .A2(net1117),
    .Y(_02344_),
    .B1(_02343_));
 sg13g2_a21oi_1 _05698_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1061),
    .A2(_02344_),
    .Y(_00050_),
    .B1(_02342_));
 sg13g2_nor2_1 _05699_ (.A(net1982),
    .B(net1059),
    .Y(_02345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05700_ (.A(net1117),
    .B_N(net1920),
    .Y(_02346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05701_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1619_[1] ),
    .A2(net1117),
    .Y(_02347_),
    .B1(_02346_));
 sg13g2_a21oi_1 _05702_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1059),
    .A2(_02347_),
    .Y(_00051_),
    .B1(_02345_));
 sg13g2_nor2b_1 _05703_ (.A(net1115),
    .B_N(\i_exotiny._1924_[26] ),
    .Y(_02348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05704_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1619_[2] ),
    .A2(net1114),
    .Y(_02349_),
    .B1(_02348_));
 sg13g2_nor2_1 _05705_ (.A(net1924),
    .B(net1058),
    .Y(_02350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05706_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1058),
    .A2(_02349_),
    .Y(_00052_),
    .B1(_02350_));
 sg13g2_nor2_1 _05707_ (.A(net1918),
    .B(net1058),
    .Y(_02351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05708_ (.A(net1115),
    .B_N(\i_exotiny._1924_[27] ),
    .Y(_02352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05709_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1619_[3] ),
    .A2(net1115),
    .Y(_02353_),
    .B1(_02352_));
 sg13g2_a21oi_1 _05710_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1058),
    .A2(_02353_),
    .Y(_00053_),
    .B1(_02351_));
 sg13g2_nor2b_1 _05711_ (.A(net1114),
    .B_N(\i_exotiny._1924_[28] ),
    .Y(_02354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05712_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1618_[0] ),
    .A2(net1114),
    .Y(_02355_),
    .B1(_02354_));
 sg13g2_nor2_1 _05713_ (.A(net1899),
    .B(net1059),
    .Y(_02356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05714_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1059),
    .A2(_02355_),
    .Y(_00054_),
    .B1(_02356_));
 sg13g2_nor2_1 _05715_ (.A(net1998),
    .B(net1059),
    .Y(_02357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05716_ (.A(net1114),
    .B_N(net1899),
    .Y(_02358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05717_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1618_[1] ),
    .A2(net1114),
    .Y(_02359_),
    .B1(_02358_));
 sg13g2_a21oi_1 _05718_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1059),
    .A2(_02359_),
    .Y(_00055_),
    .B1(_02357_));
 sg13g2_nor2_1 _05719_ (.A(net1959),
    .B(net1058),
    .Y(_02360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05720_ (.A(net1114),
    .B_N(\i_exotiny._1924_[30] ),
    .Y(_02361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05721_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1618_[2] ),
    .A2(net1114),
    .Y(_02362_),
    .B1(_02361_));
 sg13g2_a21oi_1 _05722_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1058),
    .A2(_02362_),
    .Y(_00056_),
    .B1(_02360_));
 sg13g2_nor2b_1 _05723_ (.A(net1114),
    .B_N(\i_exotiny._1924_[31] ),
    .Y(_02363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05724_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1618_[3] ),
    .A2(net1115),
    .Y(_02364_),
    .B1(_02363_));
 sg13g2_nor2_1 _05725_ (.A(net1928),
    .B(net1058),
    .Y(_02365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05726_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1058),
    .A2(_02364_),
    .Y(_00057_),
    .B1(_02365_));
 sg13g2_nand2b_1 _05727_ (.Y(_02366_),
    .B(net1105),
    .A_N(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _05728_ (.A2(_02366_),
    .A1(net2033),
    .B1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set [0]),
    .X(_00058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _05729_ (.A(\i_exotiny._1956_ ),
    .B(\i_exotiny.i_wb_spi.cnt_hbit_r[1] ),
    .C(\i_exotiny.i_wb_spi.cnt_hbit_r[2] ),
    .D(net1991),
    .Y(_02367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _05730_ (.Y(_02368_),
    .B(_02367_),
    .A_N(\i_exotiny.i_wb_spi.cnt_hbit_r[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05731_ (.Y(_02369_),
    .A(net1972),
    .B(net1073),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _05732_ (.Y(_02370_),
    .A(net1972),
    .B(_02367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05733_ (.A0(_02370_),
    .A1(\i_exotiny.i_wb_regs.spi_size_o[0] ),
    .S(net1118),
    .X(_02371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05734_ (.B1(_02369_),
    .VDD(VPWR),
    .Y(_00059_),
    .VSS(VGND),
    .A1(net1073),
    .A2(_02371_));
 sg13g2_nand2_1 _05735_ (.Y(_02372_),
    .A(\i_exotiny.i_wb_regs.spi_size_o[0] ),
    .B(\i_exotiny.i_wb_regs.spi_size_o[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _05736_ (.A(net1118),
    .B(_02372_),
    .X(_02373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05737_ (.Y(_02374_),
    .A(net1118),
    .B(_02372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05738_ (.B1(_02373_),
    .VDD(VPWR),
    .Y(_02375_),
    .VSS(VGND),
    .A1(\i_exotiny.i_wb_regs.spi_size_o[0] ),
    .A2(\i_exotiny.i_wb_regs.spi_size_o[1] ));
 sg13g2_nor2_1 _05739_ (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[5] ),
    .B(_02368_),
    .Y(_02376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _05740_ (.B(_02368_),
    .A(net3703),
    .X(_02377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05741_ (.B1(_02375_),
    .VDD(VPWR),
    .Y(_02378_),
    .VSS(VGND),
    .A1(net1118),
    .A2(_02377_));
 sg13g2_mux2_1 _05742_ (.A0(_02378_),
    .A1(net3703),
    .S(net1073),
    .X(_00060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05743_ (.A(_02373_),
    .B(_02376_),
    .Y(_02379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05744_ (.B1(net1930),
    .VDD(VPWR),
    .Y(_02380_),
    .VSS(VGND),
    .A1(_01584_),
    .A2(_02379_));
 sg13g2_nor3_1 _05745_ (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[5] ),
    .B(net1930),
    .C(_02368_),
    .Y(_02381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05746_ (.B1(_02374_),
    .VDD(VPWR),
    .Y(_02382_),
    .VSS(VGND),
    .A1(net1118),
    .A2(_02381_));
 sg13g2_o21ai_1 _05747_ (.B1(net1931),
    .VDD(VPWR),
    .Y(_00061_),
    .VSS(VGND),
    .A1(net1073),
    .A2(_02382_));
 sg13g2_and2_1 _05748_ (.A(net3606),
    .B(_01584_),
    .X(_02383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05749_ (.A(net3606),
    .B(_01584_),
    .Y(_02384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _05750_ (.A2(_02384_),
    .A1(net3634),
    .B1(_02383_),
    .X(_00062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _05751_ (.A(\i_exotiny._1956_ ),
    .B(\i_exotiny.i_wb_spi.cnt_hbit_r[1] ),
    .C(net1072),
    .Y(_02385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _05752_ (.Y(_02386_),
    .A(net3636),
    .B(_02384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05753_ (.A(_01580_),
    .B(_02386_),
    .Y(_00063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _05754_ (.Y(_02387_),
    .B(net3399),
    .A_N(_02385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _05755_ (.Y(_02388_),
    .B(_02385_),
    .A_N(net3399),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05756_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3400),
    .A2(_02388_),
    .Y(_00064_),
    .B1(_01580_));
 sg13g2_a22oi_1 _05757_ (.Y(_02389_),
    .B1(_02388_),
    .B2(net1991),
    .A2(_02367_),
    .A1(_01577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05758_ (.A(_01580_),
    .B(net1992),
    .Y(_00065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _05759_ (.Y(_02390_),
    .A(\i_exotiny._0315_[2] ),
    .B(_01465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05760_ (.Y(_02391_),
    .A(\i_exotiny._2034_[0] ),
    .B(net1127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05761_ (.Y(_02392_),
    .B1(net1126),
    .B2(net3326),
    .A2(net1144),
    .A1(net3735),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05762_ (.B1(_02392_),
    .VDD(VPWR),
    .Y(_00066_),
    .VSS(VGND),
    .A1(net1143),
    .A2(_02391_));
 sg13g2_nor3_1 _05763_ (.A(_01399_),
    .B(net1144),
    .C(net1143),
    .Y(_02393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _05764_ (.A2(net1144),
    .A1(net3553),
    .B1(_02393_),
    .X(_00067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05765_ (.Y(_02394_),
    .A(\i_exotiny._2034_[2] ),
    .B(net1127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05766_ (.Y(_02395_),
    .B1(net1126),
    .B2(net2087),
    .A2(net1144),
    .A1(net3666),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05767_ (.B1(_02395_),
    .VDD(VPWR),
    .Y(_00068_),
    .VSS(VGND),
    .A1(net1143),
    .A2(_02394_));
 sg13g2_nand2_1 _05768_ (.Y(_02396_),
    .A(\i_exotiny._2034_[3] ),
    .B(net1127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05769_ (.Y(_02397_),
    .B1(net1126),
    .B2(net2033),
    .A2(net1144),
    .A1(net3528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05770_ (.B1(_02397_),
    .VDD(VPWR),
    .Y(_00069_),
    .VSS(VGND),
    .A1(net1143),
    .A2(_02396_));
 sg13g2_nand2_1 _05771_ (.Y(_02398_),
    .A(\i_exotiny._2034_[4] ),
    .B(_00026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05772_ (.Y(_02399_),
    .B1(net1126),
    .B2(_01377_),
    .A2(net1144),
    .A1(net3785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05773_ (.B1(_02399_),
    .VDD(VPWR),
    .Y(_00070_),
    .VSS(VGND),
    .A1(net1143),
    .A2(_02398_));
 sg13g2_nand2_1 _05774_ (.Y(_02400_),
    .A(\i_exotiny._2034_[5] ),
    .B(_00026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05775_ (.Y(_02401_),
    .B1(net1126),
    .B2(_01376_),
    .A2(net1145),
    .A1(net3795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05776_ (.B1(net3796),
    .VDD(VPWR),
    .Y(_00071_),
    .VSS(VGND),
    .A1(net1143),
    .A2(_02400_));
 sg13g2_nand2_1 _05777_ (.Y(_02402_),
    .A(\i_exotiny._2034_[6] ),
    .B(net1127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05778_ (.Y(_02403_),
    .B1(net1126),
    .B2(_01375_),
    .A2(net1145),
    .A1(net3751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05779_ (.B1(net3752),
    .VDD(VPWR),
    .Y(_00072_),
    .VSS(VGND),
    .A1(net1143),
    .A2(_02402_));
 sg13g2_nand2_1 _05780_ (.Y(_02404_),
    .A(\i_exotiny._2034_[7] ),
    .B(net1127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05781_ (.Y(_02405_),
    .B1(net1126),
    .B2(_01374_),
    .A2(net1145),
    .A1(net3714),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05782_ (.B1(net3715),
    .VDD(VPWR),
    .Y(_00073_),
    .VSS(VGND),
    .A1(net1143),
    .A2(_02404_));
 sg13g2_nand2_1 _05783_ (.Y(_02406_),
    .A(\i_exotiny._2034_[8] ),
    .B(net1127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05784_ (.Y(_02407_),
    .B1(net1126),
    .B2(_01373_),
    .A2(net1145),
    .A1(net3708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05785_ (.B1(net3709),
    .VDD(VPWR),
    .Y(_00074_),
    .VSS(VGND),
    .A1(_02390_),
    .A2(_02406_));
 sg13g2_nand2_1 _05786_ (.Y(_02408_),
    .A(\i_exotiny._2034_[9] ),
    .B(_00026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05787_ (.Y(_02409_),
    .B1(_01550_),
    .B2(_01372_),
    .A2(_01549_),
    .A1(net3791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05788_ (.B1(net3792),
    .VDD(VPWR),
    .Y(_00075_),
    .VSS(VGND),
    .A1(_02390_),
    .A2(_02408_));
 sg13g2_nand2_1 _05789_ (.Y(_02410_),
    .A(\i_exotiny.i_wdg_top.o_wb_dat[10] ),
    .B(net1144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05790_ (.B1(_02410_),
    .VDD(VPWR),
    .Y(_00076_),
    .VSS(VGND),
    .A1(net1888),
    .A2(_01551_));
 sg13g2_nand2_1 _05791_ (.Y(_02411_),
    .A(net1870),
    .B(net1145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05792_ (.B1(_02411_),
    .VDD(VPWR),
    .Y(_00077_),
    .VSS(VGND),
    .A1(_00021_),
    .A2(_01551_));
 sg13g2_nand2_1 _05793_ (.Y(_02412_),
    .A(net1875),
    .B(net1145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05794_ (.B1(_02412_),
    .VDD(VPWR),
    .Y(_00078_),
    .VSS(VGND),
    .A1(_00022_),
    .A2(_01551_));
 sg13g2_nand2_1 _05795_ (.Y(_02413_),
    .A(net1873),
    .B(net1145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05796_ (.B1(_02413_),
    .VDD(VPWR),
    .Y(_00079_),
    .VSS(VGND),
    .A1(_00023_),
    .A2(_01551_));
 sg13g2_a21oi_2 _05797_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_01598_),
    .Y(_02414_),
    .A2(_01472_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_hlt_pc_ccx ));
 sg13g2_a21o_1 _05798_ (.A2(_01472_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_hlt_pc_ccx ),
    .B1(_01598_),
    .X(_02415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05799_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01605_),
    .C1(_01421_),
    .B1(_01533_),
    .A1(_01431_),
    .Y(_02416_),
    .A2(_01433_));
 sg13g2_nand4_1 _05800_ (.B(_01473_),
    .C(_01683_),
    .A(_01467_),
    .Y(_02417_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02416_));
 sg13g2_and2_1 _05801_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0] ),
    .B(_02417_),
    .X(_02418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _05802_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ),
    .C(_02418_),
    .A(net1262),
    .Y(_02419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _05803_ (.Y(_02420_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ));
 sg13g2_nor2_2 _05804_ (.A(_02419_),
    .B(_02420_),
    .Y(_02421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05805_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01443_),
    .A2(net1157),
    .Y(_02422_),
    .B1(_01473_));
 sg13g2_o21ai_1 _05806_ (.B1(net1184),
    .VDD(VPWR),
    .Y(_02423_),
    .VSS(VGND),
    .A1(\i_exotiny._1265_ ),
    .A2(net1162));
 sg13g2_a21oi_2 _05807_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_02414_),
    .Y(_02424_),
    .A2(net1142),
    .A1(_02421_));
 sg13g2_mux2_1 _05808_ (.A0(net2484),
    .A1(\i_exotiny._0018_[0] ),
    .S(net1056),
    .X(_00080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05809_ (.A0(net2815),
    .A1(\i_exotiny._0018_[1] ),
    .S(net1056),
    .X(_00081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05810_ (.A0(net2802),
    .A1(net3282),
    .S(net1056),
    .X(_00082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05811_ (.A0(net2214),
    .A1(\i_exotiny._0018_[3] ),
    .S(net1056),
    .X(_00083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05812_ (.A0(net2085),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[4] ),
    .S(net1055),
    .X(_00084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05813_ (.A0(net2321),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[5] ),
    .S(net1056),
    .X(_00085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05814_ (.A0(net2598),
    .A1(net2802),
    .S(net1057),
    .X(_00086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05815_ (.A0(net2540),
    .A1(net2214),
    .S(net1053),
    .X(_00087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05816_ (.A0(net2282),
    .A1(net2085),
    .S(net1053),
    .X(_00088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05817_ (.A0(net2750),
    .A1(net2321),
    .S(net1056),
    .X(_00089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05818_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[14] ),
    .A1(net2598),
    .S(net1057),
    .X(_00090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05819_ (.A0(net2597),
    .A1(net2540),
    .S(net1054),
    .X(_00091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05820_ (.A0(net2152),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[12] ),
    .S(net1053),
    .X(_00092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05821_ (.A0(net2745),
    .A1(net2750),
    .S(net1056),
    .X(_00093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05822_ (.A0(net2247),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[14] ),
    .S(net1057),
    .X(_00094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05823_ (.A0(net2501),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[15] ),
    .S(net1054),
    .X(_00095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05824_ (.A0(net2453),
    .A1(net2152),
    .S(net1053),
    .X(_00096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05825_ (.A0(net2543),
    .A1(net2745),
    .S(net1057),
    .X(_00097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05826_ (.A0(net2504),
    .A1(net2247),
    .S(net1054),
    .X(_00098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05827_ (.A0(net2287),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[19] ),
    .S(net1054),
    .X(_00099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05828_ (.A0(net2948),
    .A1(net2453),
    .S(net1053),
    .X(_00100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05829_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[25] ),
    .A1(net2543),
    .S(net1057),
    .X(_00101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05830_ (.A0(net2666),
    .A1(net2504),
    .S(net1054),
    .X(_00102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05831_ (.A0(net2732),
    .A1(net2287),
    .S(net1054),
    .X(_00103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05832_ (.A0(net3306),
    .A1(net2948),
    .S(net1053),
    .X(_00104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05833_ (.A0(net3370),
    .A1(net3468),
    .S(net1057),
    .X(_00105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05834_ (.A0(net2891),
    .A1(net2666),
    .S(net1054),
    .X(_00106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05835_ (.A0(net2091),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[27] ),
    .S(net1054),
    .X(_00107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05836_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1242),
    .A2(_01458_),
    .Y(_02425_),
    .B1(_01817_));
 sg13g2_a22oi_1 _05837_ (.Y(_02426_),
    .B1(_01497_),
    .B2(net1224),
    .A2(_01431_),
    .A1(_01427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05838_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1243),
    .A2(_01605_),
    .Y(_02427_),
    .B1(_01816_));
 sg13g2_and4_1 _05839_ (.A(_01610_),
    .B(_02425_),
    .C(_02426_),
    .D(_02427_),
    .X(_02428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _05840_ (.B(_02425_),
    .C(_02426_),
    .A(_01610_),
    .Y(_02429_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02427_));
 sg13g2_nand2_1 _05841_ (.Y(_02430_),
    .A(_01497_),
    .B(_02048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _05842_ (.A(_01496_),
    .B(_01497_),
    .Y(_02431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05843_ (.Y(_02432_),
    .B1(_02431_),
    .B2(_02050_),
    .A2(_02051_),
    .A1(_01496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _05844_ (.A2(_02432_),
    .A1(_02430_),
    .B1(_02429_),
    .X(_02433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _05845_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_02434_),
    .B(_02265_),
    .A(_02051_));
 sg13g2_a21oi_1 _05846_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02051_),
    .A2(_02265_),
    .Y(_02435_),
    .B1(_02428_));
 sg13g2_a21oi_1 _05847_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02434_),
    .A2(_02435_),
    .Y(_02436_),
    .B1(net1184));
 sg13g2_a22oi_1 _05848_ (.Y(_02437_),
    .B1(_02433_),
    .B2(_02436_),
    .A2(net1184),
    .A1(_01418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _05849_ (.Y(_02438_),
    .B(_02437_),
    .A_N(_01470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05850_ (.A(_02425_),
    .B_N(net1245),
    .Y(_02439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05851_ (.B1(_02439_),
    .VDD(VPWR),
    .Y(_02440_),
    .VSS(VGND),
    .A1(_02055_),
    .A2(_02069_));
 sg13g2_or3_1 _05852_ (.A(_02055_),
    .B(_02069_),
    .C(_02439_),
    .X(_02441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05853_ (.Y(_02442_),
    .A(_02440_),
    .B(_02441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05854_ (.Y(_02443_),
    .A(\i_exotiny._0352_ ),
    .B(_01470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05855_ (.B1(_02438_),
    .VDD(VPWR),
    .Y(_02444_),
    .VSS(VGND),
    .A1(_02442_),
    .A2(_02443_));
 sg13g2_mux2_1 _05856_ (.A0(net3411),
    .A1(net886),
    .S(_02421_),
    .X(_02445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05857_ (.A0(_02445_),
    .A1(net3306),
    .S(net1053),
    .X(_00108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05858_ (.B1(_02429_),
    .VDD(VPWR),
    .Y(_02446_),
    .VSS(VGND),
    .A1(_01980_),
    .A2(_02266_));
 sg13g2_a21oi_1 _05859_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01980_),
    .A2(_02266_),
    .Y(_02447_),
    .B1(_02446_));
 sg13g2_nand3_1 _05860_ (.B(_01978_),
    .C(_01979_),
    .A(_01496_),
    .Y(_02448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05861_ (.A(_01498_),
    .B(_01978_),
    .Y(_02449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05862_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01979_),
    .A2(_02431_),
    .Y(_02450_),
    .B1(_02449_));
 sg13g2_a21oi_1 _05863_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02448_),
    .A2(_02450_),
    .Y(_02451_),
    .B1(_02429_));
 sg13g2_or3_1 _05864_ (.A(net1184),
    .B(_02447_),
    .C(_02451_),
    .X(_02452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05865_ (.B1(_02452_),
    .VDD(VPWR),
    .Y(_02453_),
    .VSS(VGND),
    .A1(net3),
    .A2(_01473_));
 sg13g2_nor2_2 _05866_ (.A(_01470_),
    .B(_02453_),
    .Y(_02454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05867_ (.A0(\i_exotiny._0018_[1] ),
    .A1(net885),
    .S(_02421_),
    .X(_02455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05868_ (.A0(_02455_),
    .A1(net3370),
    .S(net1056),
    .X(_00109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05869_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01911_),
    .A2(_02267_),
    .Y(_02456_),
    .B1(_02428_));
 sg13g2_o21ai_1 _05870_ (.B1(_02456_),
    .VDD(VPWR),
    .Y(_02457_),
    .VSS(VGND),
    .A1(_01911_),
    .A2(_02267_));
 sg13g2_nor2_1 _05871_ (.A(_01498_),
    .B(_01910_),
    .Y(_02458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _05872_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01908_),
    .C1(_02458_),
    .B1(_02431_),
    .A1(_01496_),
    .Y(_02459_),
    .A2(_01911_));
 sg13g2_nor2_1 _05873_ (.A(_02429_),
    .B(_02459_),
    .Y(_02460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _05874_ (.A(net1184),
    .B(_02460_),
    .Y(_02461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _05875_ (.Y(_02462_),
    .B1(_02457_),
    .B2(_02461_),
    .A2(net1184),
    .A1(_01419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _05876_ (.A(_01470_),
    .B_N(_02462_),
    .Y(_02463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05877_ (.A0(net3282),
    .A1(net876),
    .S(_02421_),
    .X(_02464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05878_ (.A0(_02464_),
    .A1(net2891),
    .S(net1055),
    .X(_00110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _05879_ (.A(net5),
    .B(_01473_),
    .Y(_02465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _05880_ (.Y(_02466_),
    .A(_01837_),
    .B(_02268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _05881_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01836_),
    .A2(_02269_),
    .Y(_02467_),
    .B1(_02428_));
 sg13g2_a22oi_1 _05882_ (.Y(_02468_),
    .B1(_02431_),
    .B2(_01835_),
    .A2(_01836_),
    .A1(_01496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _05883_ (.B1(_02468_),
    .VDD(VPWR),
    .Y(_02469_),
    .VSS(VGND),
    .A1(_01498_),
    .A2(_01834_));
 sg13g2_a221oi_1 _05884_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02428_),
    .C1(net1184),
    .B1(_02469_),
    .A1(_02466_),
    .Y(_02470_),
    .A2(_02467_));
 sg13g2_nor2_2 _05885_ (.A(_02465_),
    .B(_02470_),
    .Y(_02471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _05886_ (.A(_01470_),
    .B(_02465_),
    .C(_02470_),
    .Y(_02472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05887_ (.A0(net2639),
    .A1(net872),
    .S(_02421_),
    .X(_02473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05888_ (.A0(_02473_),
    .A1(net2091),
    .S(net1053),
    .X(_00111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05889_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0] ),
    .B_N(_02417_),
    .Y(_02474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _05890_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ),
    .B_N(_02474_),
    .Y(_02475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _05891_ (.A(net1262),
    .B_N(_02475_),
    .Y(_02476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _05892_ (.Y(_02477_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ));
 sg13g2_nand3b_1 _05893_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .C(_02476_),
    .Y(_02478_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ));
 sg13g2_o21ai_1 _05894_ (.B1(net1158),
    .VDD(VPWR),
    .Y(_02479_),
    .VSS(VGND),
    .A1(_02423_),
    .A2(_02478_));
 sg13g2_mux2_1 _05895_ (.A0(\i_exotiny._0019_[0] ),
    .A1(net2482),
    .S(net975),
    .X(_00112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05896_ (.A0(\i_exotiny._0019_[1] ),
    .A1(net2128),
    .S(net977),
    .X(_00113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05897_ (.A0(\i_exotiny._0019_[2] ),
    .A1(net2867),
    .S(net976),
    .X(_00114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05898_ (.A0(\i_exotiny._0019_[3] ),
    .A1(net2895),
    .S(net977),
    .X(_00115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05899_ (.A0(net2482),
    .A1(net3092),
    .S(net975),
    .X(_00116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05900_ (.A0(net2128),
    .A1(net2552),
    .S(net972),
    .X(_00117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05901_ (.A0(net2867),
    .A1(net2817),
    .S(net975),
    .X(_00118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05902_ (.A0(net2895),
    .A1(net3219),
    .S(net972),
    .X(_00119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05903_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[8] ),
    .A1(net2931),
    .S(net975),
    .X(_00120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05904_ (.A0(net2552),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[13] ),
    .S(net972),
    .X(_00121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05905_ (.A0(net2817),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[14] ),
    .S(net973),
    .X(_00122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05906_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[11] ),
    .A1(net2903),
    .S(net973),
    .X(_00123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05907_ (.A0(net2931),
    .A1(net3392),
    .S(net975),
    .X(_00124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05908_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[13] ),
    .A1(net2883),
    .S(net972),
    .X(_00125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05909_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[14] ),
    .A1(net2351),
    .S(net974),
    .X(_00126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05910_ (.A0(net2903),
    .A1(net2975),
    .S(net973),
    .X(_00127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05911_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[16] ),
    .A1(net2357),
    .S(net976),
    .X(_00128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05912_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[17] ),
    .A1(net2489),
    .S(net972),
    .X(_00129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05913_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[18] ),
    .A1(net2123),
    .S(net974),
    .X(_00130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05914_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[19] ),
    .A1(net2433),
    .S(net973),
    .X(_00131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05915_ (.A0(net2357),
    .A1(net2693),
    .S(net975),
    .X(_00132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05916_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[21] ),
    .A1(net2164),
    .S(net972),
    .X(_00133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05917_ (.A0(net2123),
    .A1(net2481),
    .S(net974),
    .X(_00134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05918_ (.A0(net2433),
    .A1(net2668),
    .S(net973),
    .X(_00135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05919_ (.A0(net2693),
    .A1(net3120),
    .S(net975),
    .X(_00136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05920_ (.A0(net2164),
    .A1(net2444),
    .S(net972),
    .X(_00137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05921_ (.A0(net2481),
    .A1(net2509),
    .S(net974),
    .X(_00138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05922_ (.A0(net2668),
    .A1(net2430),
    .S(net973),
    .X(_00139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05923_ (.A0(net886),
    .A1(\i_exotiny._0019_[0] ),
    .S(_02478_),
    .X(_02480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05924_ (.A0(net3120),
    .A1(_02480_),
    .S(net975),
    .X(_00140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05925_ (.A0(net881),
    .A1(\i_exotiny._0019_[1] ),
    .S(_02478_),
    .X(_02481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05926_ (.A0(net2444),
    .A1(_02481_),
    .S(net972),
    .X(_00141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05927_ (.A0(net876),
    .A1(\i_exotiny._0019_[2] ),
    .S(_02478_),
    .X(_02482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05928_ (.A0(net2509),
    .A1(_02482_),
    .S(net973),
    .X(_00142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05929_ (.A0(net872),
    .A1(\i_exotiny._0019_[3] ),
    .S(_02478_),
    .X(_02483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05930_ (.A0(net2430),
    .A1(_02483_),
    .S(net973),
    .X(_00143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _05931_ (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ),
    .B_N(_02418_),
    .Y(_02484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _05932_ (.Y(_02485_),
    .B(_02484_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1262));
 sg13g2_nor2_2 _05933_ (.A(_02477_),
    .B(_02485_),
    .Y(_02486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _05934_ (.A2(_02486_),
    .A1(net1139),
    .B1(net1167),
    .X(_02487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05935_ (.A0(\i_exotiny._0020_[0] ),
    .A1(net2675),
    .S(net968),
    .X(_00144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05936_ (.A0(\i_exotiny._0020_[1] ),
    .A1(net3029),
    .S(net969),
    .X(_00145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05937_ (.A0(\i_exotiny._0020_[2] ),
    .A1(net2168),
    .S(net966),
    .X(_00146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05938_ (.A0(\i_exotiny._0020_[3] ),
    .A1(net3081),
    .S(net966),
    .X(_00147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05939_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[4] ),
    .A1(net2319),
    .S(net968),
    .X(_00148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05940_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[5] ),
    .A1(net2418),
    .S(net969),
    .X(_00149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05941_ (.A0(net2168),
    .A1(net3295),
    .S(net966),
    .X(_00150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05942_ (.A0(net3081),
    .A1(net3378),
    .S(net966),
    .X(_00151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05943_ (.A0(net2319),
    .A1(net2792),
    .S(net968),
    .X(_00152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05944_ (.A0(net2418),
    .A1(net3460),
    .S(net969),
    .X(_00153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05945_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[10] ),
    .A1(net2969),
    .S(net967),
    .X(_00154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05946_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[11] ),
    .A1(net2822),
    .S(net969),
    .X(_00155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05947_ (.A0(net2792),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[16] ),
    .S(net968),
    .X(_00156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05948_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[13] ),
    .A1(net2170),
    .S(net969),
    .X(_00157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05949_ (.A0(net2969),
    .A1(net3122),
    .S(net967),
    .X(_00158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05950_ (.A0(net2822),
    .A1(net2892),
    .S(net969),
    .X(_00159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05951_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[16] ),
    .A1(net3283),
    .S(net970),
    .X(_00160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05952_ (.A0(net2170),
    .A1(net3424),
    .S(net970),
    .X(_00161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05953_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[18] ),
    .A1(net2406),
    .S(net967),
    .X(_00162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05954_ (.A0(net2892),
    .A1(net2456),
    .S(net969),
    .X(_00163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05955_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[20] ),
    .A1(net2234),
    .S(net968),
    .X(_00164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05956_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[21] ),
    .A1(net2458),
    .S(net970),
    .X(_00165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05957_ (.A0(net2406),
    .A1(net2729),
    .S(net967),
    .X(_00166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05958_ (.A0(net2456),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[27] ),
    .S(net969),
    .X(_00167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05959_ (.A0(net2234),
    .A1(net2812),
    .S(net968),
    .X(_00168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05960_ (.A0(net2458),
    .A1(net2772),
    .S(net968),
    .X(_00169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05961_ (.A0(net2729),
    .A1(net2477),
    .S(net966),
    .X(_00170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05962_ (.A0(net2726),
    .A1(net2505),
    .S(net966),
    .X(_00171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05963_ (.A0(\i_exotiny._0020_[0] ),
    .A1(net888),
    .S(_02486_),
    .X(_02488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05964_ (.A0(net2812),
    .A1(_02488_),
    .S(net968),
    .X(_00172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05965_ (.A0(\i_exotiny._0020_[1] ),
    .A1(net884),
    .S(_02486_),
    .X(_02489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05966_ (.A0(net2772),
    .A1(_02489_),
    .S(net966),
    .X(_00173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05967_ (.A0(\i_exotiny._0020_[2] ),
    .A1(net878),
    .S(_02486_),
    .X(_02490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05968_ (.A0(net2477),
    .A1(_02490_),
    .S(net967),
    .X(_00174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05969_ (.A0(\i_exotiny._0020_[3] ),
    .A1(net874),
    .S(_02486_),
    .X(_02491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05970_ (.A0(net2505),
    .A1(_02491_),
    .S(net966),
    .X(_00175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _05971_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ),
    .C(_02474_),
    .Y(_02492_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1262));
 sg13g2_nor2_2 _05972_ (.A(_02420_),
    .B(_02492_),
    .Y(_02493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _05973_ (.A2(_02493_),
    .A1(net1139),
    .B1(net1167),
    .X(_02494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05974_ (.A0(\i_exotiny._0013_[0] ),
    .A1(net3417),
    .S(net1051),
    .X(_00176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05975_ (.A0(net2946),
    .A1(net3532),
    .S(net1049),
    .X(_00177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05976_ (.A0(\i_exotiny._0013_[2] ),
    .A1(net2207),
    .S(net1049),
    .X(_00178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05977_ (.A0(net2758),
    .A1(net3410),
    .S(net1051),
    .X(_00179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05978_ (.A0(net3417),
    .A1(net3484),
    .S(net1052),
    .X(_00180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05979_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[5] ),
    .A1(net2586),
    .S(net1051),
    .X(_00181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05980_ (.A0(net2207),
    .A1(net2893),
    .S(net1048),
    .X(_00182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05981_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[7] ),
    .A1(net2440),
    .S(net1051),
    .X(_00183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05982_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[8] ),
    .A1(net2154),
    .S(net1050),
    .X(_00184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05983_ (.A0(net2586),
    .A1(net2595),
    .S(net1050),
    .X(_00185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05984_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[10] ),
    .A1(net2377),
    .S(net1048),
    .X(_00186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05985_ (.A0(net2440),
    .A1(net2486),
    .S(net1051),
    .X(_00187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05986_ (.A0(net2154),
    .A1(net3234),
    .S(net1050),
    .X(_00188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05987_ (.A0(net2595),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[17] ),
    .S(net1050),
    .X(_00189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05988_ (.A0(net2377),
    .A1(net3296),
    .S(net1048),
    .X(_00190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05989_ (.A0(net2486),
    .A1(net2395),
    .S(net1051),
    .X(_00191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05990_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[16] ),
    .A1(net2343),
    .S(net1050),
    .X(_00192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05991_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[17] ),
    .A1(net3487),
    .S(net1050),
    .X(_00193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05992_ (.A0(net3296),
    .A1(net3313),
    .S(net1049),
    .X(_00194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05993_ (.A0(net2395),
    .A1(net2337),
    .S(net1051),
    .X(_00195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05994_ (.A0(net2343),
    .A1(net2754),
    .S(net1050),
    .X(_00196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05995_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[21] ),
    .A1(net2669),
    .S(net1049),
    .X(_00197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05996_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[22] ),
    .A1(net3264),
    .S(net1048),
    .X(_00198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05997_ (.A0(net2337),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[27] ),
    .S(net1051),
    .X(_00199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05998_ (.A0(net2754),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[28] ),
    .S(net1050),
    .X(_00200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _05999_ (.A0(net2669),
    .A1(net2898),
    .S(net1048),
    .X(_00201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06000_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[26] ),
    .A1(net2156),
    .S(net1048),
    .X(_00202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06001_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[27] ),
    .A1(net2630),
    .S(net1049),
    .X(_00203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06002_ (.A0(\i_exotiny._0013_[0] ),
    .A1(net887),
    .S(_02493_),
    .X(_02495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06003_ (.A0(net3513),
    .A1(_02495_),
    .S(net1049),
    .X(_00204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06004_ (.A0(net2946),
    .A1(net882),
    .S(_02493_),
    .X(_02496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06005_ (.A0(net2898),
    .A1(_02496_),
    .S(net1048),
    .X(_00205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06006_ (.A0(net2982),
    .A1(net877),
    .S(_02493_),
    .X(_02497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06007_ (.A0(net2156),
    .A1(_02497_),
    .S(net1048),
    .X(_00206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06008_ (.A0(net2758),
    .A1(net873),
    .S(_02493_),
    .X(_02498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06009_ (.A0(net2630),
    .A1(_02498_),
    .S(net1049),
    .X(_00207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06010_ (.A(_00015_),
    .B(net1105),
    .Y(_02499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06011_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3142),
    .A2(net1105),
    .Y(_00208_),
    .B1(_02499_));
 sg13g2_nor2_1 _06012_ (.A(_00016_),
    .B(net1106),
    .Y(_02500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06013_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1980),
    .A2(net1106),
    .Y(_00209_),
    .B1(_02500_));
 sg13g2_nor2_1 _06014_ (.A(_00017_),
    .B(net1106),
    .Y(_02501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06015_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2331),
    .A2(net1106),
    .Y(_00210_),
    .B1(_02501_));
 sg13g2_nor3_1 _06016_ (.A(_01465_),
    .B(_01551_),
    .C(_02126_),
    .Y(_02502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06017_ (.A(_00018_),
    .B(net1103),
    .Y(_02503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06018_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2042),
    .A2(net1103),
    .Y(_00211_),
    .B1(_02503_));
 sg13g2_nor2_1 _06019_ (.A(_00019_),
    .B(net1103),
    .Y(_02504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06020_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3559),
    .A2(net1103),
    .Y(_00212_),
    .B1(_02504_));
 sg13g2_nor2_1 _06021_ (.A(net1888),
    .B(net1104),
    .Y(_02505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06022_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3622),
    .A2(net1104),
    .Y(_00213_),
    .B1(_02505_));
 sg13g2_nor2_1 _06023_ (.A(net3543),
    .B(net1103),
    .Y(_02506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06024_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1615_[3] ),
    .A2(net1103),
    .Y(_00214_),
    .B1(_02506_));
 sg13g2_nor2_1 _06025_ (.A(_00022_),
    .B(net1103),
    .Y(_02507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06026_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2063),
    .A2(net1103),
    .Y(_00215_),
    .B1(_02507_));
 sg13g2_nor2_1 _06027_ (.A(_00023_),
    .B(net1104),
    .Y(_02508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06028_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2012),
    .A2(net1104),
    .Y(_00216_),
    .B1(_02508_));
 sg13g2_nand2_2 _06029_ (.Y(_02509_),
    .A(net1262),
    .B(_02484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06030_ (.A(_02477_),
    .B(_02509_),
    .Y(_02510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06031_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1138),
    .A2(_02510_),
    .Y(_02511_),
    .B1(net1165));
 sg13g2_mux2_1 _06032_ (.A0(net2637),
    .A1(\i_exotiny._0025_[0] ),
    .S(net964),
    .X(_00217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06033_ (.A0(net3485),
    .A1(\i_exotiny._0025_[1] ),
    .S(net963),
    .X(_00218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06034_ (.A0(net2562),
    .A1(net2521),
    .S(net962),
    .X(_00219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06035_ (.A0(net2513),
    .A1(\i_exotiny._0025_[3] ),
    .S(net963),
    .X(_00220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06036_ (.A0(net2464),
    .A1(net2637),
    .S(net964),
    .X(_00221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06037_ (.A0(net3500),
    .A1(net3485),
    .S(net962),
    .X(_00222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06038_ (.A0(net2766),
    .A1(net2562),
    .S(net962),
    .X(_00223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06039_ (.A0(net2611),
    .A1(net2513),
    .S(net963),
    .X(_00224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06040_ (.A0(net2240),
    .A1(net2464),
    .S(net964),
    .X(_00225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06041_ (.A0(net2604),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[9] ),
    .S(net961),
    .X(_00226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06042_ (.A0(net2563),
    .A1(net2766),
    .S(net962),
    .X(_00227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06043_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[15] ),
    .A1(net2611),
    .S(net963),
    .X(_00228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06044_ (.A0(net2220),
    .A1(net2240),
    .S(net961),
    .X(_00229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06045_ (.A0(net2953),
    .A1(net2604),
    .S(net961),
    .X(_00230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06046_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[18] ),
    .A1(net2563),
    .S(net962),
    .X(_00231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06047_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[19] ),
    .A1(net3060),
    .S(net963),
    .X(_00232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06048_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[20] ),
    .A1(net2220),
    .S(net965),
    .X(_00233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06049_ (.A0(net2391),
    .A1(net2953),
    .S(net961),
    .X(_00234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06050_ (.A0(net2699),
    .A1(net3025),
    .S(net961),
    .X(_00235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06051_ (.A0(net2018),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[19] ),
    .S(net964),
    .X(_00236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06052_ (.A0(net2257),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[20] ),
    .S(net964),
    .X(_00237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06053_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[25] ),
    .A1(net2391),
    .S(net961),
    .X(_00238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06054_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[26] ),
    .A1(net2699),
    .S(net961),
    .X(_00239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06055_ (.A0(net2657),
    .A1(net2018),
    .S(net963),
    .X(_00240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06056_ (.A0(net2588),
    .A1(net2257),
    .S(net964),
    .X(_00241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06057_ (.A0(net2795),
    .A1(net3389),
    .S(net961),
    .X(_00242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06058_ (.A0(net2271),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[26] ),
    .S(net962),
    .X(_00243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06059_ (.A0(net2800),
    .A1(net2657),
    .S(net963),
    .X(_00244_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06060_ (.A0(\i_exotiny._0025_[0] ),
    .A1(net887),
    .S(_02510_),
    .X(_02512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06061_ (.A0(_02512_),
    .A1(net2588),
    .S(net964),
    .X(_00245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06062_ (.A0(\i_exotiny._0025_[1] ),
    .A1(net882),
    .S(_02510_),
    .X(_02513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06063_ (.A0(_02513_),
    .A1(net2795),
    .S(net962),
    .X(_00246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06064_ (.A0(net2521),
    .A1(net877),
    .S(_02510_),
    .X(_02514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06065_ (.A0(_02514_),
    .A1(net2271),
    .S(net962),
    .X(_00247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06066_ (.A0(\i_exotiny._0025_[3] ),
    .A1(net873),
    .S(_02510_),
    .X(_02515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06067_ (.A0(_02515_),
    .A1(net2800),
    .S(net963),
    .X(_00248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06068_ (.Y(_02516_),
    .A(net2140),
    .B(_01701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06069_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01739_),
    .A2(_02516_),
    .Y(_00249_),
    .B1(_01388_));
 sg13g2_nand2_2 _06070_ (.Y(_02517_),
    .A(net1262),
    .B(_02475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _06071_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_02518_),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ));
 sg13g2_nor2_2 _06072_ (.A(_02517_),
    .B(_02518_),
    .Y(_02519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _06073_ (.A2(_02519_),
    .A1(net1139),
    .B1(net1166),
    .X(_02520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06074_ (.A0(net2933),
    .A1(net3461),
    .S(net957),
    .X(_00250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06075_ (.A0(net2791),
    .A1(net3091),
    .S(net956),
    .X(_00251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06076_ (.A0(\i_exotiny._0038_[2] ),
    .A1(net2255),
    .S(net959),
    .X(_00252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06077_ (.A0(\i_exotiny._0038_[3] ),
    .A1(net2303),
    .S(net960),
    .X(_00253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06078_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[4] ),
    .A1(net3349),
    .S(net957),
    .X(_00254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06079_ (.A0(net3091),
    .A1(net3193),
    .S(net955),
    .X(_00255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06080_ (.A0(net2255),
    .A1(net2843),
    .S(net958),
    .X(_00256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06081_ (.A0(net2303),
    .A1(net2761),
    .S(net960),
    .X(_00257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06082_ (.A0(net3349),
    .A1(net3423),
    .S(net955),
    .X(_00258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06083_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[9] ),
    .A1(net2148),
    .S(net955),
    .X(_00259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06084_ (.A0(net2843),
    .A1(net3131),
    .S(net958),
    .X(_00260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06085_ (.A0(net2761),
    .A1(net3366),
    .S(net960),
    .X(_00261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06086_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[12] ),
    .A1(net2844),
    .S(net956),
    .X(_00262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06087_ (.A0(net2148),
    .A1(net3316),
    .S(net955),
    .X(_00263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06088_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[14] ),
    .A1(net2619),
    .S(net958),
    .X(_00264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06089_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[15] ),
    .A1(net2073),
    .S(net960),
    .X(_00265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06090_ (.A0(net2844),
    .A1(net3428),
    .S(net956),
    .X(_00266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06091_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[17] ),
    .A1(net3279),
    .S(net955),
    .X(_00267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06092_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[18] ),
    .A1(net2413),
    .S(net958),
    .X(_00268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06093_ (.A0(net2073),
    .A1(net2855),
    .S(net960),
    .X(_00269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06094_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[20] ),
    .A1(net2798),
    .S(net956),
    .X(_00270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06095_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[21] ),
    .A1(net2593),
    .S(net955),
    .X(_00271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06096_ (.A0(net2413),
    .A1(net2769),
    .S(net958),
    .X(_00272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06097_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[23] ),
    .A1(net2435),
    .S(net958),
    .X(_00273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06098_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[24] ),
    .A1(net2276),
    .S(net957),
    .X(_00274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06099_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[25] ),
    .A1(net2400),
    .S(net955),
    .X(_00275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06100_ (.A0(net2769),
    .A1(net2756),
    .S(net958),
    .X(_00276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06101_ (.A0(net2435),
    .A1(net3169),
    .S(net959),
    .X(_00277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06102_ (.A0(net2933),
    .A1(net888),
    .S(_02519_),
    .X(_02521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06103_ (.A0(net2276),
    .A1(_02521_),
    .S(net957),
    .X(_00278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06104_ (.A0(net2791),
    .A1(net883),
    .S(_02519_),
    .X(_02522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06105_ (.A0(net2400),
    .A1(_02522_),
    .S(net955),
    .X(_00279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06106_ (.A0(\i_exotiny._0038_[2] ),
    .A1(net878),
    .S(_02519_),
    .X(_02523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06107_ (.A0(net2756),
    .A1(_02523_),
    .S(net958),
    .X(_00280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06108_ (.A0(net3412),
    .A1(net874),
    .S(_02519_),
    .X(_02524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06109_ (.A0(net3169),
    .A1(_02524_),
    .S(net959),
    .X(_00281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _06110_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ),
    .C(_02418_),
    .Y(_02525_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1262));
 sg13g2_nor2_2 _06111_ (.A(_02518_),
    .B(_02525_),
    .Y(_02526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _06112_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net1165),
    .Y(_02527_),
    .A2(_02526_),
    .A1(net1138));
 sg13g2_mux2_1 _06113_ (.A0(net3111),
    .A1(\i_exotiny._0037_[0] ),
    .S(net1043),
    .X(_00282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06114_ (.A0(net2317),
    .A1(\i_exotiny._0037_[1] ),
    .S(net1047),
    .X(_00283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06115_ (.A0(net2961),
    .A1(\i_exotiny._0037_[2] ),
    .S(net1047),
    .X(_00284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06116_ (.A0(net2115),
    .A1(\i_exotiny._0037_[3] ),
    .S(net1046),
    .X(_00285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06117_ (.A0(net2762),
    .A1(net3111),
    .S(net1043),
    .X(_00286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06118_ (.A0(net2539),
    .A1(net2317),
    .S(net1047),
    .X(_00287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06119_ (.A0(net2691),
    .A1(net2961),
    .S(net1047),
    .X(_00288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06120_ (.A0(net2632),
    .A1(net2115),
    .S(net1046),
    .X(_00289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06121_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[12] ),
    .A1(net2762),
    .S(net1043),
    .X(_00290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06122_ (.A0(net2979),
    .A1(net2539),
    .S(net1046),
    .X(_00291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06123_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[14] ),
    .A1(net2691),
    .S(net1045),
    .X(_00292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06124_ (.A0(net2602),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[11] ),
    .S(net1044),
    .X(_00293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06125_ (.A0(net3014),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[12] ),
    .S(net1043),
    .X(_00294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06126_ (.A0(net3038),
    .A1(net2979),
    .S(net1046),
    .X(_00295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06127_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[18] ),
    .A1(net3450),
    .S(net1045),
    .X(_00296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06128_ (.A0(net3454),
    .A1(net2602),
    .S(net1044),
    .X(_00297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06129_ (.A0(net3005),
    .A1(net3014),
    .S(net1043),
    .X(_00298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06130_ (.A0(net3171),
    .A1(net3038),
    .S(net1047),
    .X(_00299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06131_ (.A0(net2261),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[18] ),
    .S(net1045),
    .X(_00300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06132_ (.A0(net3503),
    .A1(net3454),
    .S(net1044),
    .X(_00301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06133_ (.A0(net2709),
    .A1(net3005),
    .S(net1043),
    .X(_00302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06134_ (.A0(net2389),
    .A1(net3171),
    .S(net1047),
    .X(_00303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06135_ (.A0(net3011),
    .A1(net2261),
    .S(net1045),
    .X(_00304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06136_ (.A0(net2333),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[23] ),
    .S(net1044),
    .X(_00305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06137_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[28] ),
    .A1(net2709),
    .S(net1043),
    .X(_00306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06138_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[29] ),
    .A1(net2389),
    .S(net1046),
    .X(_00307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06139_ (.A0(net2664),
    .A1(net3011),
    .S(net1045),
    .X(_00308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06140_ (.A0(net2658),
    .A1(net2333),
    .S(net1046),
    .X(_00309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06141_ (.A0(\i_exotiny._0037_[0] ),
    .A1(net887),
    .S(_02526_),
    .X(_02528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06142_ (.A0(_02528_),
    .A1(net3302),
    .S(net1043),
    .X(_00310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06143_ (.A0(\i_exotiny._0037_[1] ),
    .A1(net882),
    .S(_02526_),
    .X(_02529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06144_ (.A0(_02529_),
    .A1(net2682),
    .S(net1046),
    .X(_00311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06145_ (.A0(\i_exotiny._0037_[2] ),
    .A1(net877),
    .S(_02526_),
    .X(_02530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06146_ (.A0(_02530_),
    .A1(net2664),
    .S(net1045),
    .X(_00312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06147_ (.A0(net3442),
    .A1(net873),
    .S(_02526_),
    .X(_02531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06148_ (.A0(_02531_),
    .A1(net2658),
    .S(net1046),
    .X(_00313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _06149_ (.Y(_02532_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ),
    .B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _06150_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .C(_02476_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ),
    .Y(_02533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06151_ (.B1(net1158),
    .VDD(VPWR),
    .Y(_02534_),
    .VSS(VGND),
    .A1(_02423_),
    .A2(_02533_));
 sg13g2_mux2_1 _06152_ (.A0(\i_exotiny._0028_[0] ),
    .A1(net3127),
    .S(net953),
    .X(_00314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06153_ (.A0(\i_exotiny._0028_[1] ),
    .A1(net3393),
    .S(net951),
    .X(_00315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06154_ (.A0(\i_exotiny._0028_[2] ),
    .A1(net2166),
    .S(net952),
    .X(_00316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06155_ (.A0(\i_exotiny._0028_[3] ),
    .A1(net3102),
    .S(net950),
    .X(_00317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06156_ (.A0(net3127),
    .A1(net3191),
    .S(net954),
    .X(_00318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06157_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[5] ),
    .A1(net3277),
    .S(net951),
    .X(_00319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06158_ (.A0(net2166),
    .A1(net2557),
    .S(net952),
    .X(_00320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06159_ (.A0(net3102),
    .A1(net2739),
    .S(net950),
    .X(_00321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06160_ (.A0(net3191),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[12] ),
    .S(net953),
    .X(_00322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06161_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[9] ),
    .A1(net2218),
    .S(net953),
    .X(_00323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06162_ (.A0(net2557),
    .A1(net3149),
    .S(net952),
    .X(_00324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06163_ (.A0(net2739),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[15] ),
    .S(net950),
    .X(_00325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06164_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[12] ),
    .A1(net3245),
    .S(net954),
    .X(_00326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06165_ (.A0(net2218),
    .A1(net2873),
    .S(net952),
    .X(_00327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06166_ (.A0(net3149),
    .A1(net3441),
    .S(net952),
    .X(_00328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06167_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[15] ),
    .A1(net2263),
    .S(net950),
    .X(_00329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06168_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[16] ),
    .A1(net2109),
    .S(net953),
    .X(_00330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06169_ (.A0(net2873),
    .A1(net3096),
    .S(net951),
    .X(_00331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06170_ (.A0(net3441),
    .A1(net3435),
    .S(net952),
    .X(_00332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06171_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[19] ),
    .A1(net2238),
    .S(net950),
    .X(_00333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06172_ (.A0(net2109),
    .A1(net2554),
    .S(net953),
    .X(_00334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06173_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[21] ),
    .A1(net2226),
    .S(net951),
    .X(_00335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06174_ (.A0(net3435),
    .A1(net3398),
    .S(net953),
    .X(_00336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06175_ (.A0(net2238),
    .A1(net2591),
    .S(net950),
    .X(_00337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06176_ (.A0(net2554),
    .A1(net2768),
    .S(net953),
    .X(_00338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06177_ (.A0(net2226),
    .A1(net3023),
    .S(net951),
    .X(_00339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06178_ (.A0(net3398),
    .A1(net3161),
    .S(net952),
    .X(_00340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06179_ (.A0(net2591),
    .A1(net3174),
    .S(net950),
    .X(_00341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06180_ (.A0(net890),
    .A1(net3269),
    .S(_02533_),
    .X(_02535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06181_ (.A0(net2768),
    .A1(_02535_),
    .S(net954),
    .X(_00342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06182_ (.A0(net885),
    .A1(\i_exotiny._0028_[1] ),
    .S(_02533_),
    .X(_02536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06183_ (.A0(net3023),
    .A1(_02536_),
    .S(net951),
    .X(_00343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06184_ (.A0(net876),
    .A1(\i_exotiny._0028_[2] ),
    .S(_02533_),
    .X(_02537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06185_ (.A0(net3161),
    .A1(_02537_),
    .S(net952),
    .X(_00344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06186_ (.A0(_02472_),
    .A1(net3212),
    .S(_02533_),
    .X(_02538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06187_ (.A0(net3174),
    .A1(_02538_),
    .S(net950),
    .X(_00345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06188_ (.Y(_02539_),
    .A(_01365_),
    .B(net1105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06189_ (.A2(_02539_),
    .A1(net2087),
    .B1(net1263),
    .X(_00346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06190_ (.A(_02509_),
    .B(_02532_),
    .Y(_02540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06191_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1140),
    .A2(_02540_),
    .Y(_02541_),
    .B1(net1166));
 sg13g2_mux2_1 _06192_ (.A0(net2146),
    .A1(\i_exotiny._0033_[0] ),
    .S(net948),
    .X(_00347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06193_ (.A0(net2230),
    .A1(\i_exotiny._0033_[1] ),
    .S(net945),
    .X(_00348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06194_ (.A0(net2565),
    .A1(net3337),
    .S(net948),
    .X(_00349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06195_ (.A0(net3495),
    .A1(net3510),
    .S(net946),
    .X(_00350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06196_ (.A0(net2629),
    .A1(net2146),
    .S(net948),
    .X(_00351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06197_ (.A0(net2947),
    .A1(net2230),
    .S(net945),
    .X(_00352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06198_ (.A0(net2427),
    .A1(net2565),
    .S(net948),
    .X(_00353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06199_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[11] ),
    .A1(net3495),
    .S(net947),
    .X(_00354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06200_ (.A0(net3205),
    .A1(net2629),
    .S(net947),
    .X(_00355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06201_ (.A0(net3186),
    .A1(net2947),
    .S(net946),
    .X(_00356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06202_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[14] ),
    .A1(net2427),
    .S(net948),
    .X(_00357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06203_ (.A0(net3479),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[11] ),
    .S(net949),
    .X(_00358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06204_ (.A0(net2863),
    .A1(net3205),
    .S(net947),
    .X(_00359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06205_ (.A0(net2643),
    .A1(net3186),
    .S(net946),
    .X(_00360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06206_ (.A0(net2566),
    .A1(net2794),
    .S(net948),
    .X(_00361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06207_ (.A0(net3188),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[15] ),
    .S(net947),
    .X(_00362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06208_ (.A0(net2375),
    .A1(net2863),
    .S(net947),
    .X(_00363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06209_ (.A0(net2369),
    .A1(net2643),
    .S(net946),
    .X(_00364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06210_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[22] ),
    .A1(net2566),
    .S(net948),
    .X(_00365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06211_ (.A0(net2475),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[19] ),
    .S(net949),
    .X(_00366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06212_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[24] ),
    .A1(net2375),
    .S(net947),
    .X(_00367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06213_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[25] ),
    .A1(net2369),
    .S(net946),
    .X(_00368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06214_ (.A0(net2774),
    .A1(net3427),
    .S(net945),
    .X(_00369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06215_ (.A0(net2717),
    .A1(net2475),
    .S(net947),
    .X(_00370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06216_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[28] ),
    .A1(net2479),
    .S(net948),
    .X(_00371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06217_ (.A0(net2305),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[25] ),
    .S(net945),
    .X(_00372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06218_ (.A0(net2671),
    .A1(net2774),
    .S(net945),
    .X(_00373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06219_ (.A0(net3208),
    .A1(net2717),
    .S(net947),
    .X(_00374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06220_ (.A0(\i_exotiny._0033_[0] ),
    .A1(net888),
    .S(_02540_),
    .X(_02542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06221_ (.A0(_02542_),
    .A1(net3455),
    .S(net945),
    .X(_00375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06222_ (.A0(net2871),
    .A1(net883),
    .S(_02540_),
    .X(_02543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06223_ (.A0(_02543_),
    .A1(net2305),
    .S(net945),
    .X(_00376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06224_ (.A0(\i_exotiny._0033_[2] ),
    .A1(net878),
    .S(_02540_),
    .X(_02544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06225_ (.A0(_02544_),
    .A1(net2671),
    .S(net945),
    .X(_00377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06226_ (.A0(\i_exotiny._0033_[3] ),
    .A1(net874),
    .S(_02540_),
    .X(_02545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06227_ (.A0(_02545_),
    .A1(net3208),
    .S(net946),
    .X(_00378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06228_ (.A(_02525_),
    .B(_02532_),
    .Y(_02546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06229_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1139),
    .A2(_02546_),
    .Y(_02547_),
    .B1(net1166));
 sg13g2_mux2_1 _06230_ (.A0(net2095),
    .A1(\i_exotiny._0031_[0] ),
    .S(net1040),
    .X(_00379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06231_ (.A0(net3515),
    .A1(\i_exotiny._0031_[1] ),
    .S(net1040),
    .X(_00380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06232_ (.A0(net3336),
    .A1(net3231),
    .S(net1041),
    .X(_00381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06233_ (.A0(net2136),
    .A1(\i_exotiny._0031_[3] ),
    .S(net1039),
    .X(_00382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06234_ (.A0(net2986),
    .A1(net2095),
    .S(net1040),
    .X(_00383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06235_ (.A0(net2416),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[5] ),
    .S(net1040),
    .X(_00384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06236_ (.A0(net3087),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[6] ),
    .S(net1038),
    .X(_00385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06237_ (.A0(net2415),
    .A1(net2136),
    .S(net1039),
    .X(_00386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06238_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[12] ),
    .A1(net2986),
    .S(net1040),
    .X(_00387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06239_ (.A0(net3211),
    .A1(net2416),
    .S(net1040),
    .X(_00388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06240_ (.A0(net3334),
    .A1(net3087),
    .S(net1038),
    .X(_00389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06241_ (.A0(net2914),
    .A1(net2415),
    .S(net1039),
    .X(_00390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06242_ (.A0(net2621),
    .A1(net3213),
    .S(net1041),
    .X(_00391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06243_ (.A0(net2894),
    .A1(net3211),
    .S(net1041),
    .X(_00392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06244_ (.A0(net3285),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[14] ),
    .S(net1038),
    .X(_00393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06245_ (.A0(net2939),
    .A1(net2914),
    .S(net1039),
    .X(_00394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06246_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[20] ),
    .A1(net2621),
    .S(net1041),
    .X(_00395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06247_ (.A0(net2373),
    .A1(net2894),
    .S(net1041),
    .X(_00396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06248_ (.A0(net2180),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[18] ),
    .S(net1038),
    .X(_00397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06249_ (.A0(net3357),
    .A1(net2939),
    .S(net1038),
    .X(_00398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06250_ (.A0(net2200),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[20] ),
    .S(net1041),
    .X(_00399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06251_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[25] ),
    .A1(net2373),
    .S(net1040),
    .X(_00400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06252_ (.A0(net2915),
    .A1(net2180),
    .S(net1038),
    .X(_00401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06253_ (.A0(net3159),
    .A1(net3357),
    .S(net1038),
    .X(_00402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06254_ (.A0(net2741),
    .A1(net2200),
    .S(net1041),
    .X(_00403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06255_ (.A0(net3164),
    .A1(net3409),
    .S(net1039),
    .X(_00404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06256_ (.A0(net3136),
    .A1(net2915),
    .S(net1038),
    .X(_00405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06257_ (.A0(net2640),
    .A1(net3159),
    .S(net1039),
    .X(_00406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06258_ (.A0(net3123),
    .A1(net888),
    .S(_02546_),
    .X(_02548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06259_ (.A0(_02548_),
    .A1(net2741),
    .S(net1040),
    .X(_00407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06260_ (.A0(\i_exotiny._0031_[1] ),
    .A1(net883),
    .S(_02546_),
    .X(_02549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06261_ (.A0(_02549_),
    .A1(net3164),
    .S(net1039),
    .X(_00408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06262_ (.A0(net3231),
    .A1(net878),
    .S(_02546_),
    .X(_02550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06263_ (.A0(_02550_),
    .A1(net3136),
    .S(net1042),
    .X(_00409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06264_ (.A0(\i_exotiny._0031_[3] ),
    .A1(net874),
    .S(_02546_),
    .X(_02551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06265_ (.A0(_02551_),
    .A1(net2640),
    .S(net1039),
    .X(_00410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06266_ (.A(_02420_),
    .B(_02509_),
    .Y(_02552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06267_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1140),
    .A2(_02552_),
    .Y(_02553_),
    .B1(net1166));
 sg13g2_mux2_1 _06268_ (.A0(net3179),
    .A1(\i_exotiny._0016_[0] ),
    .S(net942),
    .X(_00411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06269_ (.A0(net2119),
    .A1(\i_exotiny._0016_[1] ),
    .S(net939),
    .X(_00412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06270_ (.A0(net3026),
    .A1(\i_exotiny._0016_[2] ),
    .S(net939),
    .X(_00413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06271_ (.A0(net2647),
    .A1(net2814),
    .S(net943),
    .X(_00414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06272_ (.A0(net2402),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[4] ),
    .S(net942),
    .X(_00415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06273_ (.A0(net2881),
    .A1(net2119),
    .S(net939),
    .X(_00416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06274_ (.A0(net3348),
    .A1(net3026),
    .S(net939),
    .X(_00417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06275_ (.A0(net2385),
    .A1(net2647),
    .S(net943),
    .X(_00418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06276_ (.A0(net2708),
    .A1(net2402),
    .S(net942),
    .X(_00419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06277_ (.A0(net2832),
    .A1(net2881),
    .S(net939),
    .X(_00420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06278_ (.A0(net2775),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[10] ),
    .S(net941),
    .X(_00421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06279_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[15] ),
    .A1(net2385),
    .S(net942),
    .X(_00422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06280_ (.A0(net2507),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[12] ),
    .S(net942),
    .X(_00423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06281_ (.A0(net2797),
    .A1(net2832),
    .S(net940),
    .X(_00424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06282_ (.A0(net2963),
    .A1(net2775),
    .S(net944),
    .X(_00425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06283_ (.A0(net3405),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[15] ),
    .S(net943),
    .X(_00426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06284_ (.A0(net2698),
    .A1(net2507),
    .S(net942),
    .X(_00427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06285_ (.A0(net2367),
    .A1(net2797),
    .S(net940),
    .X(_00428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06286_ (.A0(net3332),
    .A1(net2963),
    .S(net941),
    .X(_00429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06287_ (.A0(net2820),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[19] ),
    .S(net943),
    .X(_00430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06288_ (.A0(net2778),
    .A1(net2698),
    .S(net941),
    .X(_00431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06289_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[25] ),
    .A1(net2367),
    .S(net940),
    .X(_00432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06290_ (.A0(net3229),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[22] ),
    .S(net941),
    .X(_00433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06291_ (.A0(net2887),
    .A1(net2820),
    .S(net943),
    .X(_00434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06292_ (.A0(net2383),
    .A1(net2778),
    .S(net941),
    .X(_00435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06293_ (.A0(net2424),
    .A1(net3362),
    .S(net940),
    .X(_00436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06294_ (.A0(net3206),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[26] ),
    .S(net939),
    .X(_00437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06295_ (.A0(net2673),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[27] ),
    .S(net942),
    .X(_00438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06296_ (.A0(\i_exotiny._0016_[0] ),
    .A1(net888),
    .S(_02552_),
    .X(_02554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06297_ (.A0(_02554_),
    .A1(net2383),
    .S(net941),
    .X(_00439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06298_ (.A0(\i_exotiny._0016_[1] ),
    .A1(net884),
    .S(_02552_),
    .X(_02555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06299_ (.A0(_02555_),
    .A1(net2424),
    .S(net939),
    .X(_00440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06300_ (.A0(net3274),
    .A1(net878),
    .S(_02552_),
    .X(_02556_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06301_ (.A0(_02556_),
    .A1(net3206),
    .S(net939),
    .X(_00441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06302_ (.A0(net2814),
    .A1(net875),
    .S(_02552_),
    .X(_02557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06303_ (.A0(_02557_),
    .A1(net2673),
    .S(net942),
    .X(_00442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06304_ (.A(_02420_),
    .B(_02525_),
    .Y(_02558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06305_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1138),
    .A2(_02558_),
    .Y(_02559_),
    .B1(net1165));
 sg13g2_mux2_1 _06306_ (.A0(net3429),
    .A1(net3260),
    .S(net1034),
    .X(_00443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06307_ (.A0(net2465),
    .A1(\i_exotiny._0014_[1] ),
    .S(net1033),
    .X(_00444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06308_ (.A0(net3519),
    .A1(net3674),
    .S(net1037),
    .X(_00445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06309_ (.A0(net3263),
    .A1(net3044),
    .S(net1033),
    .X(_00446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06310_ (.A0(net2426),
    .A1(net3429),
    .S(net1035),
    .X(_00447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06311_ (.A0(net2538),
    .A1(net2465),
    .S(net1033),
    .X(_00448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06312_ (.A0(net3478),
    .A1(net3519),
    .S(net1036),
    .X(_00449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06313_ (.A0(net2826),
    .A1(net3263),
    .S(net1033),
    .X(_00450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06314_ (.A0(net2325),
    .A1(net2426),
    .S(net1036),
    .X(_00451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06315_ (.A0(net2650),
    .A1(net2538),
    .S(net1034),
    .X(_00452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06316_ (.A0(net3257),
    .A1(net3478),
    .S(net1036),
    .X(_00453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06317_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[15] ),
    .A1(net2826),
    .S(net1033),
    .X(_00454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06318_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[16] ),
    .A1(net2325),
    .S(net1035),
    .X(_00455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06319_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[17] ),
    .A1(net2650),
    .S(net1034),
    .X(_00456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06320_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[18] ),
    .A1(net3257),
    .S(net1036),
    .X(_00457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06321_ (.A0(net3266),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[15] ),
    .S(net1036),
    .X(_00458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06322_ (.A0(net1976),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[16] ),
    .S(net1035),
    .X(_00459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06323_ (.A0(net2113),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[17] ),
    .S(net1034),
    .X(_00460_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06324_ (.A0(net2949),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[18] ),
    .S(net1035),
    .X(_00461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06325_ (.A0(net2000),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[19] ),
    .S(net1036),
    .X(_00462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06326_ (.A0(net2429),
    .A1(net1976),
    .S(net1035),
    .X(_00463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06327_ (.A0(net2730),
    .A1(net2113),
    .S(net1034),
    .X(_00464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06328_ (.A0(net2016),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[22] ),
    .S(net1035),
    .X(_00465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06329_ (.A0(net2719),
    .A1(net2000),
    .S(net1033),
    .X(_00466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06330_ (.A0(net3223),
    .A1(net2429),
    .S(net1035),
    .X(_00467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06331_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[29] ),
    .A1(net2730),
    .S(net1034),
    .X(_00468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06332_ (.A0(net2353),
    .A1(net2016),
    .S(net1035),
    .X(_00469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06333_ (.A0(net2971),
    .A1(net2719),
    .S(net1037),
    .X(_00470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06334_ (.A0(net3260),
    .A1(net887),
    .S(_02558_),
    .X(_02560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06335_ (.A0(_02560_),
    .A1(net3223),
    .S(net1034),
    .X(_00471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06336_ (.A0(\i_exotiny._0014_[1] ),
    .A1(net882),
    .S(_02558_),
    .X(_02561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06337_ (.A0(_02561_),
    .A1(net3147),
    .S(net1033),
    .X(_00472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06338_ (.A0(\i_exotiny._0014_[2] ),
    .A1(net877),
    .S(_02558_),
    .X(_02562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06339_ (.A0(_02562_),
    .A1(net2353),
    .S(net1036),
    .X(_00473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06340_ (.A0(net3044),
    .A1(net873),
    .S(_02558_),
    .X(_02563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06341_ (.A0(_02563_),
    .A1(net2971),
    .S(net1033),
    .X(_00474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _06342_ (.B(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ),
    .C(_02474_),
    .A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ),
    .Y(_02564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06343_ (.A(_02532_),
    .B(_02564_),
    .Y(_02565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06344_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1140),
    .A2(_02565_),
    .Y(_02566_),
    .B1(net1167));
 sg13g2_mux2_1 _06345_ (.A0(net2138),
    .A1(\i_exotiny._0035_[0] ),
    .S(net1029),
    .X(_00475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06346_ (.A0(net3261),
    .A1(net3419),
    .S(net1029),
    .X(_00476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06347_ (.A0(net3373),
    .A1(net3343),
    .S(net1030),
    .X(_00477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06348_ (.A0(net3539),
    .A1(\i_exotiny._0035_[3] ),
    .S(net1031),
    .X(_00478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06349_ (.A0(net2929),
    .A1(net2138),
    .S(net1029),
    .X(_00479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06350_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[9] ),
    .A1(net3261),
    .S(net1028),
    .X(_00480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06351_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[10] ),
    .A1(net3373),
    .S(net1030),
    .X(_00481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06352_ (.A0(net2269),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[7] ),
    .S(net1030),
    .X(_00482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06353_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[12] ),
    .A1(net2929),
    .S(net1029),
    .X(_00483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06354_ (.A0(net3354),
    .A1(net3379),
    .S(net1028),
    .X(_00484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06355_ (.A0(net2283),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[10] ),
    .S(net1032),
    .X(_00485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06356_ (.A0(net2851),
    .A1(net2269),
    .S(net1030),
    .X(_00486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06357_ (.A0(net3432),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[12] ),
    .S(net1028),
    .X(_00487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06358_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[17] ),
    .A1(net3354),
    .S(net1028),
    .X(_00488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06359_ (.A0(net2292),
    .A1(net2283),
    .S(net1031),
    .X(_00489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06360_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[19] ),
    .A1(net2851),
    .S(net1030),
    .X(_00490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06361_ (.A0(net2493),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[16] ),
    .S(net1028),
    .X(_00491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06362_ (.A0(net2473),
    .A1(net3439),
    .S(net1031),
    .X(_00492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06363_ (.A0(net2764),
    .A1(net2292),
    .S(net1032),
    .X(_00493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06364_ (.A0(net2515),
    .A1(net2942),
    .S(net1030),
    .X(_00494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06365_ (.A0(net2995),
    .A1(net2493),
    .S(net1028),
    .X(_00495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06366_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[25] ),
    .A1(net2473),
    .S(net1031),
    .X(_00496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06367_ (.A0(net2196),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[22] ),
    .S(net1031),
    .X(_00497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06368_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[27] ),
    .A1(net2515),
    .S(net1031),
    .X(_00498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06369_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[28] ),
    .A1(net2995),
    .S(net1028),
    .X(_00499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06370_ (.A0(net2576),
    .A1(net3053),
    .S(net1028),
    .X(_00500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06371_ (.A0(net2718),
    .A1(net2196),
    .S(net1031),
    .X(_00501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06372_ (.A0(net2522),
    .A1(net3135),
    .S(net1030),
    .X(_00502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06373_ (.A0(\i_exotiny._0035_[0] ),
    .A1(net889),
    .S(_02565_),
    .X(_02567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06374_ (.A0(_02567_),
    .A1(net3324),
    .S(net1029),
    .X(_00503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06375_ (.A0(\i_exotiny._0035_[1] ),
    .A1(net884),
    .S(_02565_),
    .X(_02568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06376_ (.A0(_02568_),
    .A1(net2576),
    .S(net1029),
    .X(_00504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06377_ (.A0(net3343),
    .A1(net879),
    .S(_02565_),
    .X(_02569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06378_ (.A0(_02569_),
    .A1(net2718),
    .S(net1030),
    .X(_00505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06379_ (.A0(\i_exotiny._0035_[3] ),
    .A1(net875),
    .S(_02565_),
    .X(_02570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06380_ (.A0(_02570_),
    .A1(net2522),
    .S(net1029),
    .X(_00506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06381_ (.B1(_01513_),
    .VDD(VPWR),
    .Y(_02571_),
    .VSS(VGND),
    .A1(_01489_),
    .A2(_01521_));
 sg13g2_nand2_1 _06382_ (.Y(_02572_),
    .A(_01524_),
    .B(_02571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06383_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3702),
    .A2(net10),
    .Y(_02573_),
    .B1(net1225));
 sg13g2_nand2_1 _06384_ (.Y(_00507_),
    .A(_02572_),
    .B(_02573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _06385_ (.A(net3775),
    .B(_01484_),
    .C(_01489_),
    .D(_01521_),
    .Y(_02574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06386_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3647),
    .A2(_02180_),
    .Y(_02575_),
    .B1(_02574_));
 sg13g2_nor2_1 _06387_ (.A(net1225),
    .B(net3648),
    .Y(_00508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06388_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3764),
    .A2(_02180_),
    .Y(_02576_),
    .B1(net1225));
 sg13g2_o21ai_1 _06389_ (.B1(_02576_),
    .VDD(VPWR),
    .Y(_00509_),
    .VSS(VGND),
    .A1(_01513_),
    .A2(_02131_));
 sg13g2_nand2_1 _06390_ (.Y(_02577_),
    .A(net3493),
    .B(net1271),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06391_ (.B1(_02577_),
    .VDD(VPWR),
    .Y(_02578_),
    .VSS(VGND),
    .A1(net1273),
    .A2(_01391_));
 sg13g2_nor2_1 _06392_ (.A(_02574_),
    .B(_02578_),
    .Y(_02579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06393_ (.A(_02219_),
    .B(_02572_),
    .C(_02579_),
    .Y(_02580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06394_ (.A2(net1071),
    .A1(net3787),
    .B1(_02580_),
    .X(_00510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06395_ (.A0(\i_exotiny._0315_[8] ),
    .A1(net3476),
    .S(net1272),
    .X(_02581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _06396_ (.Y(_02582_),
    .B1(_02581_),
    .B2(_01525_),
    .A2(_02180_),
    .A1(net3828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06397_ (.Y(_00511_),
    .A(net1284),
    .B(net3829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06398_ (.A0(net3665),
    .A1(net3509),
    .S(net1272),
    .X(_02583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06399_ (.A(_02574_),
    .B(_02583_),
    .Y(_02584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06400_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3778),
    .A2(_02180_),
    .Y(_02585_),
    .B1(net1225));
 sg13g2_o21ai_1 _06401_ (.B1(_02585_),
    .VDD(VPWR),
    .Y(_00512_),
    .VSS(VGND),
    .A1(_02572_),
    .A2(_02584_));
 sg13g2_mux2_1 _06402_ (.A0(\i_exotiny._0315_[16] ),
    .A1(\i_exotiny._0314_[16] ),
    .S(net1271),
    .X(_02586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _06403_ (.Y(_02587_),
    .B1(_02586_),
    .B2(_01512_),
    .A2(_01520_),
    .A1(_01485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06404_ (.A(_01522_),
    .B(_02586_),
    .Y(_02588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06405_ (.A(_02219_),
    .B(_02587_),
    .C(_02588_),
    .Y(_02589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06406_ (.A2(net1071),
    .A1(net3759),
    .B1(_02589_),
    .X(_00513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06407_ (.Y(_02590_),
    .A(net2014),
    .B(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06408_ (.A0(\i_exotiny._0315_[20] ),
    .A1(\i_exotiny._0314_[20] ),
    .S(net1271),
    .X(_02591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _06409_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02591_),
    .C1(_01553_),
    .B1(_02571_),
    .A1(_01520_),
    .Y(_02592_),
    .A2(_02226_));
 sg13g2_o21ai_1 _06410_ (.B1(_02590_),
    .VDD(VPWR),
    .Y(_00514_),
    .VSS(VGND),
    .A1(_02219_),
    .A2(_02592_));
 sg13g2_nor3_2 _06411_ (.A(_01390_),
    .B(net1233),
    .C(\i_exotiny._0315_[4] ),
    .Y(_02593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _06412_ (.B(net1219),
    .C(net1146),
    .A(_01437_),
    .Y(_02594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _06413_ (.B(net1219),
    .C(net1146),
    .A(_01437_),
    .Y(_02595_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02593_));
 sg13g2_nand3_1 _06414_ (.B(net1146),
    .C(_02593_),
    .A(_01447_),
    .Y(_02596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06415_ (.A(\i_exotiny._0327_[0] ),
    .B(net3688),
    .C(_02596_),
    .Y(_02597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06416_ (.B1(net1282),
    .VDD(VPWR),
    .Y(_02598_),
    .VSS(VGND),
    .A1(_01361_),
    .A2(_02595_));
 sg13g2_a21o_1 _06417_ (.A2(_02595_),
    .A1(net3551),
    .B1(_02598_),
    .X(_00515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06418_ (.B1(net1282),
    .VDD(VPWR),
    .Y(_02599_),
    .VSS(VGND),
    .A1(_01366_),
    .A2(_02595_));
 sg13g2_a21o_1 _06419_ (.A2(_02595_),
    .A1(net3618),
    .B1(_02599_),
    .X(_00516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06420_ (.A(net3730),
    .B(_02595_),
    .Y(_02600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06421_ (.B1(net1282),
    .VDD(VPWR),
    .Y(_02601_),
    .VSS(VGND),
    .A1(net3561),
    .A2(net3689));
 sg13g2_nor2_1 _06422_ (.A(_02600_),
    .B(_02601_),
    .Y(_00517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06423_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3430),
    .A2(_02595_),
    .Y(_02602_),
    .B1(net1227));
 sg13g2_nand2_1 _06424_ (.Y(_02603_),
    .A(net3611),
    .B(net3689),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06425_ (.Y(_00518_),
    .A(_02602_),
    .B(_02603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06426_ (.A(_01489_),
    .B(_01513_),
    .Y(_02604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06427_ (.B1(net1284),
    .VDD(VPWR),
    .Y(_02605_),
    .VSS(VGND),
    .A1(net3775),
    .A2(_02604_));
 sg13g2_inv_1 _06428_ (.VDD(VPWR),
    .Y(_00519_),
    .A(net3776),
    .VSS(VGND));
 sg13g2_nand3_1 _06429_ (.B(net1146),
    .C(_02593_),
    .A(net1219),
    .Y(_02606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _06430_ (.A(net1225),
    .B(_02130_),
    .C(_02606_),
    .Y(_02607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06431_ (.A0(net3733),
    .A1(net3717),
    .S(_02607_),
    .X(_00520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06432_ (.A0(net3721),
    .A1(net3697),
    .S(_02607_),
    .X(_00521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06433_ (.A(_02509_),
    .B(_02518_),
    .Y(_02608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _06434_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net1165),
    .Y(_02609_),
    .A2(_02608_),
    .A1(net1138));
 sg13g2_mux2_1 _06435_ (.A0(net2905),
    .A1(\i_exotiny._0039_[0] ),
    .S(net938),
    .X(_00522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06436_ (.A0(net3037),
    .A1(net3064),
    .S(net936),
    .X(_00523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06437_ (.A0(net2777),
    .A1(net3291),
    .S(net937),
    .X(_00524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06438_ (.A0(net3344),
    .A1(\i_exotiny._0039_[3] ),
    .S(net934),
    .X(_00525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06439_ (.A0(net2609),
    .A1(net2905),
    .S(net937),
    .X(_00526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06440_ (.A0(net2232),
    .A1(net3037),
    .S(net934),
    .X(_00527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06441_ (.A0(net2550),
    .A1(net2777),
    .S(net937),
    .X(_00528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06442_ (.A0(net2057),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[7] ),
    .S(net934),
    .X(_00529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06443_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[12] ),
    .A1(net2609),
    .S(net937),
    .X(_00530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06444_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[13] ),
    .A1(net2232),
    .S(net934),
    .X(_00531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06445_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[14] ),
    .A1(net2550),
    .S(_02609_),
    .X(_00532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06446_ (.A0(net2206),
    .A1(net2057),
    .S(net935),
    .X(_00533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06447_ (.A0(net2737),
    .A1(net3003),
    .S(net937),
    .X(_00534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06448_ (.A0(net2381),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[13] ),
    .S(net934),
    .X(_00535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06449_ (.A0(net2648),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[14] ),
    .S(net938),
    .X(_00536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06450_ (.A0(net2679),
    .A1(net2206),
    .S(net935),
    .X(_00537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06451_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[20] ),
    .A1(net2737),
    .S(net938),
    .X(_00538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06452_ (.A0(net2955),
    .A1(net2381),
    .S(net934),
    .X(_00539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06453_ (.A0(net2667),
    .A1(net2648),
    .S(net938),
    .X(_00540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06454_ (.A0(net3166),
    .A1(net2679),
    .S(net935),
    .X(_00541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06455_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[24] ),
    .A1(net3068),
    .S(net938),
    .X(_00542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06456_ (.A0(net3172),
    .A1(net2955),
    .S(net934),
    .X(_00543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06457_ (.A0(net3342),
    .A1(net2667),
    .S(net937),
    .X(_00544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06458_ (.A0(net3115),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[23] ),
    .S(net935),
    .X(_00545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06459_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[28] ),
    .A1(net3151),
    .S(net938),
    .X(_00546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06460_ (.A0(net2249),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[25] ),
    .S(net934),
    .X(_00547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06461_ (.A0(net3322),
    .A1(net3342),
    .S(net937),
    .X(_00548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06462_ (.A0(net3346),
    .A1(net3115),
    .S(net935),
    .X(_00549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06463_ (.A0(\i_exotiny._0039_[0] ),
    .A1(net886),
    .S(_02608_),
    .X(_02610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06464_ (.A0(_02610_),
    .A1(net3328),
    .S(net938),
    .X(_00550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06465_ (.A0(net3064),
    .A1(net881),
    .S(_02608_),
    .X(_02611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06466_ (.A0(_02611_),
    .A1(net2249),
    .S(net936),
    .X(_00551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06467_ (.A0(net3291),
    .A1(net877),
    .S(_02608_),
    .X(_02612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06468_ (.A0(_02612_),
    .A1(net3322),
    .S(net937),
    .X(_00552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06469_ (.A0(\i_exotiny._0039_[3] ),
    .A1(net873),
    .S(_02608_),
    .X(_02613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06470_ (.A0(_02613_),
    .A1(net3346),
    .S(net935),
    .X(_00553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06471_ (.A(_02419_),
    .B(_02518_),
    .Y(_02614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _06472_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net1166),
    .Y(_02615_),
    .A2(_02614_),
    .A1(net1139));
 sg13g2_mux2_1 _06473_ (.A0(net3351),
    .A1(net2703),
    .S(net1024),
    .X(_00554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06474_ (.A0(net2983),
    .A1(net3133),
    .S(net1024),
    .X(_00555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06475_ (.A0(net3482),
    .A1(\i_exotiny._0041_[2] ),
    .S(net1025),
    .X(_00556_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06476_ (.A0(net2081),
    .A1(\i_exotiny._0041_[3] ),
    .S(net1023),
    .X(_00557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06477_ (.A0(net3297),
    .A1(net3351),
    .S(net1024),
    .X(_00558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06478_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[9] ),
    .A1(net2983),
    .S(net1025),
    .X(_00559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06479_ (.A0(net2530),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[6] ),
    .S(net1027),
    .X(_00560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06480_ (.A0(net2578),
    .A1(net2081),
    .S(net1023),
    .X(_00561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06481_ (.A0(net3022),
    .A1(net3297),
    .S(net1023),
    .X(_00562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06482_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[13] ),
    .A1(net3019),
    .S(net1025),
    .X(_00563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06483_ (.A0(net3298),
    .A1(net2530),
    .S(net1026),
    .X(_00564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06484_ (.A0(net3195),
    .A1(net2578),
    .S(net1023),
    .X(_00565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06485_ (.A0(net2448),
    .A1(net3022),
    .S(net1026),
    .X(_00566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06486_ (.A0(net2876),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[13] ),
    .S(net1025),
    .X(_00567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06487_ (.A0(net3021),
    .A1(net3298),
    .S(net1026),
    .X(_00568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06488_ (.A0(net2940),
    .A1(net3195),
    .S(net1023),
    .X(_00569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06489_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[20] ),
    .A1(net2448),
    .S(net1026),
    .X(_00570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06490_ (.A0(net3101),
    .A1(net2876),
    .S(net1025),
    .X(_00571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06491_ (.A0(net3012),
    .A1(net3021),
    .S(net1027),
    .X(_00572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06492_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[23] ),
    .A1(net2940),
    .S(net1023),
    .X(_00573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06493_ (.A0(net2228),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[20] ),
    .S(net1026),
    .X(_00574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06494_ (.A0(net2583),
    .A1(net3101),
    .S(net1027),
    .X(_00575_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06495_ (.A0(net2659),
    .A1(net3012),
    .S(net1026),
    .X(_00576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06496_ (.A0(net2363),
    .A1(net2999),
    .S(net1023),
    .X(_00577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06497_ (.A0(net2561),
    .A1(net2228),
    .S(net1026),
    .X(_00578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06498_ (.A0(net2532),
    .A1(net2583),
    .S(net1025),
    .X(_00579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06499_ (.A0(net2341),
    .A1(net2659),
    .S(net1026),
    .X(_00580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06500_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[31] ),
    .A1(net2363),
    .S(net1023),
    .X(_00581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06501_ (.A0(net2703),
    .A1(net888),
    .S(_02614_),
    .X(_02616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06502_ (.A0(_02616_),
    .A1(net2561),
    .S(net1024),
    .X(_00582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06503_ (.A0(\i_exotiny._0041_[1] ),
    .A1(net883),
    .S(_02614_),
    .X(_02617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06504_ (.A0(_02617_),
    .A1(net2532),
    .S(net1025),
    .X(_00583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06505_ (.A0(\i_exotiny._0041_[2] ),
    .A1(net878),
    .S(_02614_),
    .X(_02618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06506_ (.A0(_02618_),
    .A1(net2341),
    .S(net1025),
    .X(_00584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06507_ (.A0(\i_exotiny._0041_[3] ),
    .A1(net874),
    .S(_02614_),
    .X(_02619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06508_ (.A0(_02619_),
    .A1(net3117),
    .S(net1024),
    .X(_00585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06509_ (.A(_02420_),
    .B(_02485_),
    .Y(_02620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _06510_ (.A2(_02620_),
    .A1(net1142),
    .B1(net1160),
    .X(_02621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06511_ (.A0(net3031),
    .A1(net2835),
    .S(net932),
    .X(_00586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06512_ (.A0(\i_exotiny._0043_[1] ),
    .A1(net2285),
    .S(net932),
    .X(_00587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06513_ (.A0(\i_exotiny._0043_[2] ),
    .A1(net3094),
    .S(net930),
    .X(_00588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06514_ (.A0(\i_exotiny._0043_[3] ),
    .A1(net2274),
    .S(net931),
    .X(_00589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06515_ (.A0(net2835),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[8] ),
    .S(net932),
    .X(_00590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06516_ (.A0(net2285),
    .A1(net2541),
    .S(net932),
    .X(_00591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06517_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[6] ),
    .A1(net2824),
    .S(net929),
    .X(_00592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06518_ (.A0(net2274),
    .A1(net2590),
    .S(net930),
    .X(_00593_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06519_ (.A0(net3153),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[12] ),
    .S(net932),
    .X(_00594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06520_ (.A0(net2541),
    .A1(net3132),
    .S(net932),
    .X(_00595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06521_ (.A0(net2824),
    .A1(net2902),
    .S(net929),
    .X(_00596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06522_ (.A0(net2590),
    .A1(net2606),
    .S(net930),
    .X(_00597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06523_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[12] ),
    .A1(net2874),
    .S(net933),
    .X(_00598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06524_ (.A0(net3132),
    .A1(net3054),
    .S(net932),
    .X(_00599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06525_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[14] ),
    .A1(net2184),
    .S(net929),
    .X(_00600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06526_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[15] ),
    .A1(net2224),
    .S(net930),
    .X(_00601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06527_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[16] ),
    .A1(net2701),
    .S(net933),
    .X(_00602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06528_ (.A0(net3054),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[21] ),
    .S(net931),
    .X(_00603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06529_ (.A0(net2184),
    .A1(net2437),
    .S(net929),
    .X(_00604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06530_ (.A0(net2224),
    .A1(net2943),
    .S(net930),
    .X(_00605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06531_ (.A0(net2701),
    .A1(net2919),
    .S(net933),
    .X(_00606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06532_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[21] ),
    .A1(net2623),
    .S(net931),
    .X(_00607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06533_ (.A0(net2437),
    .A1(net2965),
    .S(net929),
    .X(_00608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06534_ (.A0(net2943),
    .A1(net2782),
    .S(net930),
    .X(_00609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06535_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[24] ),
    .A1(net2617),
    .S(net933),
    .X(_00610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06536_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[25] ),
    .A1(net2150),
    .S(net931),
    .X(_00611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06537_ (.A0(net2965),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[30] ),
    .S(net929),
    .X(_00612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06538_ (.A0(net2782),
    .A1(net2491),
    .S(net930),
    .X(_00613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06539_ (.A0(net3031),
    .A1(net886),
    .S(_02620_),
    .X(_02622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06540_ (.A0(net2617),
    .A1(_02622_),
    .S(net932),
    .X(_00614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06541_ (.A0(net2753),
    .A1(net881),
    .S(_02620_),
    .X(_02623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06542_ (.A0(net2150),
    .A1(_02623_),
    .S(net929),
    .X(_00615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06543_ (.A0(\i_exotiny._0043_[2] ),
    .A1(net876),
    .S(_02620_),
    .X(_02624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06544_ (.A0(net3239),
    .A1(_02624_),
    .S(net929),
    .X(_00616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06545_ (.A0(\i_exotiny._0043_[3] ),
    .A1(net872),
    .S(_02620_),
    .X(_02625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06546_ (.A0(net2491),
    .A1(_02625_),
    .S(net930),
    .X(_00617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06547_ (.A0(\i_exotiny._0369_[7] ),
    .A1(net3591),
    .S(net1210),
    .X(_00618_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _06548_ (.A(\i_exotiny._0369_[8] ),
    .B(net1213),
    .X(_02626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06549_ (.A2(net1210),
    .A1(net3757),
    .B1(_02626_),
    .X(_00619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06550_ (.A(net1262),
    .B(net1215),
    .Y(_02627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06551_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01406_),
    .A2(net1216),
    .Y(_00620_),
    .B1(_02627_));
 sg13g2_and2_1 _06552_ (.A(net3443),
    .B(net1213),
    .X(_02628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06553_ (.A2(net1210),
    .A1(net3794),
    .B1(_02628_),
    .X(_00621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _06554_ (.A(net3641),
    .B(net1213),
    .X(_02629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06555_ (.A2(net1210),
    .A1(net3783),
    .B1(_02629_),
    .X(_00622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06556_ (.A0(net1261),
    .A1(net3596),
    .S(net1216),
    .X(_00623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06557_ (.A0(net3787),
    .A1(net1259),
    .S(net1211),
    .X(_00624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06558_ (.A0(net3810),
    .A1(net3675),
    .S(net1216),
    .X(_00625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06559_ (.A0(net3818),
    .A1(net3737),
    .S(net1216),
    .X(_00626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06560_ (.A(net3505),
    .B(_01504_),
    .Y(_02630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06561_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01394_),
    .A2(net1211),
    .Y(_00627_),
    .B1(_02630_));
 sg13g2_nor2_1 _06562_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ),
    .B(net1160),
    .Y(_02631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06563_ (.A(net3493),
    .B(net1152),
    .Y(_02632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06564_ (.A(net1195),
    .B(_02631_),
    .C(_02632_),
    .Y(_00628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06565_ (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ),
    .B(net1160),
    .Y(_02633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06566_ (.A(net3603),
    .B(net1154),
    .Y(_02634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06567_ (.A(net1200),
    .B(_02633_),
    .C(_02634_),
    .Y(_00629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06568_ (.A(\i_exotiny._0314_[2] ),
    .B(net1162),
    .Y(_02635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06569_ (.A(net3407),
    .B(net1155),
    .Y(_02636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06570_ (.A(net1200),
    .B(_02635_),
    .C(_02636_),
    .Y(_00630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06571_ (.A(net3390),
    .B(net1162),
    .Y(_02637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06572_ (.A(net3605),
    .B(net1156),
    .Y(_02638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06573_ (.A(net1200),
    .B(_02637_),
    .C(_02638_),
    .Y(_00631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06574_ (.A(\i_exotiny._0314_[4] ),
    .B(net1160),
    .Y(_02639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06575_ (.A(net3476),
    .B(net1152),
    .Y(_02640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06576_ (.A(net1194),
    .B(_02639_),
    .C(_02640_),
    .Y(_00632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06577_ (.A(\i_exotiny._0314_[5] ),
    .B(net1162),
    .Y(_02641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06578_ (.A(net3382),
    .B(net1155),
    .Y(_02642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06579_ (.A(net1199),
    .B(_02641_),
    .C(_02642_),
    .Y(_00633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06580_ (.A(net3407),
    .B(net1164),
    .Y(_02643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06581_ (.A(net3475),
    .B(net1156),
    .Y(_02644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06582_ (.A(net1199),
    .B(_02643_),
    .C(_02644_),
    .Y(_00634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06583_ (.A(\i_exotiny._0314_[7] ),
    .B(net1164),
    .Y(_02645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06584_ (.A(net3517),
    .B(net1155),
    .Y(_02646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06585_ (.A(net1199),
    .B(_02645_),
    .C(_02646_),
    .Y(_00635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06586_ (.A(net3476),
    .B(net1159),
    .Y(_02647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06587_ (.A(net3509),
    .B(net1153),
    .Y(_02648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06588_ (.A(net1194),
    .B(_02647_),
    .C(_02648_),
    .Y(_00636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06589_ (.A(net3382),
    .B(net1162),
    .Y(_02649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06590_ (.A(net3504),
    .B(net1154),
    .Y(_02650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06591_ (.A(net1199),
    .B(_02649_),
    .C(_02650_),
    .Y(_00637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06592_ (.A(\i_exotiny._0314_[10] ),
    .B(net1163),
    .Y(_02651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06593_ (.A(net3462),
    .B(net1156),
    .Y(_02652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06594_ (.A(net1198),
    .B(_02651_),
    .C(_02652_),
    .Y(_00638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06595_ (.A(\i_exotiny._0314_[11] ),
    .B(net1163),
    .Y(_02653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06596_ (.A(net3498),
    .B(net1155),
    .Y(_02654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06597_ (.A(net1198),
    .B(_02653_),
    .C(_02654_),
    .Y(_00639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06598_ (.A(\i_exotiny._0314_[12] ),
    .B(net1159),
    .Y(_02655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06599_ (.A(net3447),
    .B(net1153),
    .Y(_02656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06600_ (.A(net1194),
    .B(_02655_),
    .C(_02656_),
    .Y(_00640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06601_ (.A(\i_exotiny._0314_[13] ),
    .B(net1160),
    .Y(_02657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06602_ (.A(net2864),
    .B(net1154),
    .Y(_02658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06603_ (.A(net1198),
    .B(_02657_),
    .C(_02658_),
    .Y(_00641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06604_ (.A(\i_exotiny._0314_[14] ),
    .B(net1163),
    .Y(_02659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06605_ (.A(net3402),
    .B(net1156),
    .Y(_02660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06606_ (.A(net1199),
    .B(_02659_),
    .C(_02660_),
    .Y(_00642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06607_ (.A(\i_exotiny._0314_[15] ),
    .B(net1163),
    .Y(_02661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06608_ (.A(net3243),
    .B(net1155),
    .Y(_02662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06609_ (.A(net1198),
    .B(_02661_),
    .C(_02662_),
    .Y(_00643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06610_ (.A(\i_exotiny._0314_[16] ),
    .B(net1159),
    .Y(_02663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06611_ (.A(net3358),
    .B(net1152),
    .Y(_02664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06612_ (.A(net1194),
    .B(_02663_),
    .C(_02664_),
    .Y(_00644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06613_ (.A(net2864),
    .B(net1160),
    .Y(_02665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06614_ (.A(net3489),
    .B(net1157),
    .Y(_02666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06615_ (.A(net1194),
    .B(_02665_),
    .C(_02666_),
    .Y(_00645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06616_ (.A(net3402),
    .B(net1163),
    .Y(_02667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06617_ (.A(net3610),
    .B(net1155),
    .Y(_02668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06618_ (.A(net1199),
    .B(_02667_),
    .C(_02668_),
    .Y(_00646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06619_ (.A(\i_exotiny._0314_[19] ),
    .B(net1160),
    .Y(_02669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06620_ (.A(net3155),
    .B(net1155),
    .Y(_02670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06621_ (.A(net1198),
    .B(_02669_),
    .C(_02670_),
    .Y(_00647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06622_ (.A(\i_exotiny._0314_[20] ),
    .B(net1159),
    .Y(_02671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06623_ (.A(net2038),
    .B(net1152),
    .Y(_02672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06624_ (.A(net1195),
    .B(_02671_),
    .C(_02672_),
    .Y(_00648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06625_ (.A(\i_exotiny._0314_[21] ),
    .B(net1159),
    .Y(_02673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06626_ (.A(net2008),
    .B(net1152),
    .Y(_02674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06627_ (.A(net1194),
    .B(_02673_),
    .C(_02674_),
    .Y(_00649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06628_ (.A(\i_exotiny._0314_[22] ),
    .B(net1161),
    .Y(_02675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06629_ (.A(net1965),
    .B(net1155),
    .Y(_02676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06630_ (.A(net1199),
    .B(_02675_),
    .C(_02676_),
    .Y(_00650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06631_ (.A(\i_exotiny._0314_[23] ),
    .B(net1161),
    .Y(_02677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06632_ (.A(net1974),
    .B(net1154),
    .Y(_02678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06633_ (.A(net1198),
    .B(_02677_),
    .C(_02678_),
    .Y(_00651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06634_ (.A(net2038),
    .B(net1159),
    .Y(_02679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06635_ (.A(net2446),
    .B(net1152),
    .Y(_02680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06636_ (.A(net1195),
    .B(_02679_),
    .C(_02680_),
    .Y(_00652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06637_ (.A(net2008),
    .B(net1159),
    .Y(_02681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06638_ (.A(net2002),
    .B(net1153),
    .Y(_02682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06639_ (.A(net1194),
    .B(_02681_),
    .C(_02682_),
    .Y(_00653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06640_ (.A(net1965),
    .B(net1161),
    .Y(_02683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06641_ (.A(net2886),
    .B(net1154),
    .Y(_02684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06642_ (.A(net1198),
    .B(_02683_),
    .C(_02684_),
    .Y(_00654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06643_ (.A(net1974),
    .B(net1161),
    .Y(_02685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06644_ (.A(net2037),
    .B(net1154),
    .Y(_02686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06645_ (.A(net1198),
    .B(_02685_),
    .C(_02686_),
    .Y(_00655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06646_ (.Y(_02687_),
    .A(net2446),
    .B(net1152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _06647_ (.A(net1268),
    .B(_01461_),
    .C(_02440_),
    .D(_02441_),
    .X(_02688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _06648_ (.B(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r [0]),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ),
    .X(_02689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06649_ (.A(_01388_),
    .B(_01467_),
    .Y(_02690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _06650_ (.Y(_02691_),
    .A(net1269),
    .B(_01466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06651_ (.A0(_02689_),
    .A1(_02437_),
    .S(_02688_),
    .X(_02692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06652_ (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data [0]),
    .B(_02691_),
    .Y(_02693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06653_ (.A(\i_exotiny._0352_ ),
    .B(net1153),
    .C(_02693_),
    .Y(_02694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06654_ (.B1(_02694_),
    .VDD(VPWR),
    .Y(_02695_),
    .VSS(VGND),
    .A1(_02690_),
    .A2(_02692_));
 sg13g2_a21oi_1 _06655_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02687_),
    .A2(_02695_),
    .Y(_00656_),
    .B1(net1195));
 sg13g2_nand2_1 _06656_ (.Y(_02696_),
    .A(net2002),
    .B(net1152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06657_ (.A2(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r [0]),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ),
    .B1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ),
    .X(_02697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06658_ (.Y(_02698_),
    .A(_02259_),
    .B(_02697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06659_ (.A0(_02698_),
    .A1(_02453_),
    .S(_02688_),
    .X(_02699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06660_ (.B1(net1162),
    .VDD(VPWR),
    .Y(_02700_),
    .VSS(VGND),
    .A1(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data [0]),
    .A2(_02691_));
 sg13g2_a21o_1 _06661_ (.A2(_02699_),
    .A1(_02691_),
    .B1(_02700_),
    .X(_02701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06662_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02696_),
    .A2(_02701_),
    .Y(_00657_),
    .B1(net1194));
 sg13g2_xnor2_1 _06663_ (.Y(_02702_),
    .A(\i_exotiny._0314_[2] ),
    .B(_02262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _06664_ (.Y(_02703_),
    .B(_02688_),
    .A_N(_02462_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06665_ (.B1(_02691_),
    .VDD(VPWR),
    .Y(_02704_),
    .VSS(VGND),
    .A1(_02688_),
    .A2(_02702_));
 sg13g2_nand2b_1 _06666_ (.Y(_02705_),
    .B(_02703_),
    .A_N(_02704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06667_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3730),
    .A2(_02690_),
    .Y(_02706_),
    .B1(net1153));
 sg13g2_a221oi_1 _06668_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02706_),
    .C1(net1196),
    .B1(_02705_),
    .A1(_01370_),
    .Y(_00658_),
    .A2(net1154));
 sg13g2_o21ai_1 _06669_ (.B1(_02688_),
    .VDD(VPWR),
    .Y(_02707_),
    .VSS(VGND),
    .A1(_02465_),
    .A2(_02470_));
 sg13g2_xor2_1 _06670_ (.B(_02263_),
    .A(net3390),
    .X(_02708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06671_ (.B1(_02691_),
    .VDD(VPWR),
    .Y(_02709_),
    .VSS(VGND),
    .A1(_02688_),
    .A2(_02708_));
 sg13g2_nand2b_1 _06672_ (.Y(_02710_),
    .B(_02707_),
    .A_N(_02709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06673_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3611),
    .A2(_02690_),
    .Y(_02711_),
    .B1(net1153));
 sg13g2_a221oi_1 _06674_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02711_),
    .C1(net1195),
    .B1(_02710_),
    .A1(_01369_),
    .Y(_00659_),
    .A2(net1153));
 sg13g2_nand4_1 _06675_ (.B(net1224),
    .C(net1234),
    .A(net1249),
    .Y(_02712_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01463_));
 sg13g2_nand4_1 _06676_ (.B(\i_exotiny._0327_[0] ),
    .C(_01464_),
    .A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ),
    .Y(_02713_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01532_));
 sg13g2_a21oi_1 _06677_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01362_),
    .A2(_02712_),
    .Y(_02714_),
    .B1(_02713_));
 sg13g2_and3_1 _06678_ (.X(_02715_),
    .A(net1270),
    .B(_01388_),
    .C(net1137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06679_ (.A(_01362_),
    .B(_02712_),
    .Y(_02716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _06680_ (.A(_02714_),
    .B(_02715_),
    .C(_02716_),
    .Y(_02717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _06681_ (.Y(_02718_),
    .A(net1102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06682_ (.A(_01506_),
    .B(_02718_),
    .Y(_02719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06683_ (.Y(_02720_),
    .A(net1137),
    .B(net1102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _06684_ (.Y(_02721_),
    .B(net1219),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1181));
 sg13g2_nor3_1 _06685_ (.A(\i_exotiny._0315_[3] ),
    .B(net1233),
    .C(_01391_),
    .Y(_02722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _06686_ (.X(_02723_),
    .A(_01390_),
    .B(net1233),
    .C(_01391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _06687_ (.Y(_02724_),
    .B1(_02723_),
    .B2(net15),
    .A2(_02593_),
    .A1(net3551),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _06688_ (.A(_02593_),
    .B(_02722_),
    .C(_02723_),
    .Y(_02725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _06689_ (.Y(_02726_),
    .B1(_02725_),
    .B2(\i_exotiny.gpo[0] ),
    .A2(_02722_),
    .A1(net1116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06690_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02724_),
    .A2(_02726_),
    .Y(_02727_),
    .B1(_02721_));
 sg13g2_nand2b_1 _06691_ (.Y(_02728_),
    .B(net1187),
    .A_N(net2014),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06692_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01407_),
    .A2(net1193),
    .Y(_02729_),
    .B1(net1169));
 sg13g2_a221oi_1 _06693_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02729_),
    .C1(_02727_),
    .B1(_02728_),
    .A1(\i_exotiny.i_wdg_top.o_wb_dat[0] ),
    .Y(_02730_),
    .A2(net1181));
 sg13g2_nor2_1 _06694_ (.A(net3632),
    .B(net1102),
    .Y(_02731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _06695_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01506_),
    .C1(_02731_),
    .B1(_02730_),
    .A1(_01361_),
    .Y(_00660_),
    .A2(_02719_));
 sg13g2_nand2_1 _06696_ (.Y(_02732_),
    .A(net3741),
    .B(_02725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06697_ (.Y(_02733_),
    .A(net3576),
    .B(net1193),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _06698_ (.Y(_02734_),
    .B1(_02723_),
    .B2(net16),
    .A2(_02593_),
    .A1(net3618),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _06699_ (.B(_02732_),
    .C(_02734_),
    .A(net1219),
    .Y(_02735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06700_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[1] ),
    .A2(net1187),
    .Y(_02736_),
    .B1(net1219));
 sg13g2_a21oi_1 _06701_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02733_),
    .A2(_02736_),
    .Y(_02737_),
    .B1(net1181));
 sg13g2_a221oi_1 _06702_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02737_),
    .C1(net1137),
    .B1(_02735_),
    .A1(net3553),
    .Y(_02738_),
    .A2(net1181));
 sg13g2_a221oi_1 _06703_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01366_),
    .C1(_02738_),
    .B1(_02719_),
    .A1(_01392_),
    .Y(_00661_),
    .A2(net1068));
 sg13g2_nand2_1 _06704_ (.Y(_02739_),
    .A(\i_exotiny.gpo[2] ),
    .B(_02725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _06705_ (.Y(_02740_),
    .B1(_02723_),
    .B2(net17),
    .A2(_02593_),
    .A1(\i_exotiny._2025_[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06706_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02739_),
    .A2(_02740_),
    .Y(_02741_),
    .B1(_02721_));
 sg13g2_mux2_1 _06707_ (.A0(\i_exotiny._0369_[2] ),
    .A1(net3574),
    .S(net1193),
    .X(_02742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _06708_ (.A(net3719),
    .B(net1102),
    .Y(_02743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _06709_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02742_),
    .C1(_02741_),
    .B1(net1173),
    .A1(net3666),
    .Y(_02744_),
    .A2(net1181));
 sg13g2_a221oi_1 _06710_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01506_),
    .C1(_02743_),
    .B1(_02744_),
    .A1(_01365_),
    .Y(_00662_),
    .A2(_02719_));
 sg13g2_nor4_2 _06711_ (.A(_01390_),
    .B(net1233),
    .C(\i_exotiny._0315_[4] ),
    .Y(_02745_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_02721_));
 sg13g2_mux2_1 _06712_ (.A0(\i_exotiny._0369_[3] ),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[3] ),
    .S(net1193),
    .X(_02746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _06713_ (.A(_02721_),
    .B_N(_02723_),
    .Y(_02747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _06714_ (.Y(_02748_),
    .B1(_02746_),
    .B2(net1173),
    .A2(_02745_),
    .A1(net3430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _06715_ (.Y(_02749_),
    .B1(_02747_),
    .B2(net6),
    .A2(net1182),
    .A1(net3528),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06716_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02748_),
    .A2(_02749_),
    .Y(_02750_),
    .B1(net1137));
 sg13g2_a21oi_1 _06717_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3611),
    .A2(net1137),
    .Y(_02751_),
    .B1(_02750_));
 sg13g2_nor2_1 _06718_ (.A(net3657),
    .B(net1102),
    .Y(_02752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06719_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1102),
    .A2(_02751_),
    .Y(_00663_),
    .B1(_02752_));
 sg13g2_o21ai_1 _06720_ (.B1(net1173),
    .VDD(VPWR),
    .Y(_02753_),
    .VSS(VGND),
    .A1(net3654),
    .A2(net1187));
 sg13g2_a21oi_1 _06721_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01403_),
    .A2(net1187),
    .Y(_02754_),
    .B1(_02753_));
 sg13g2_a221oi_1 _06722_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net7),
    .C1(_02754_),
    .B1(_02747_),
    .A1(net3785),
    .Y(_02755_),
    .A2(net1182));
 sg13g2_a22oi_1 _06723_ (.Y(_02756_),
    .B1(_02719_),
    .B2(net3808),
    .A2(net1068),
    .A1(net3567),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06724_ (.B1(_02756_),
    .VDD(VPWR),
    .Y(_00664_),
    .VSS(VGND),
    .A1(net1137),
    .A2(_02755_));
 sg13g2_nor2_1 _06725_ (.A(net3142),
    .B(_02720_),
    .Y(_02757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06726_ (.B1(net1173),
    .VDD(VPWR),
    .Y(_02758_),
    .VSS(VGND),
    .A1(\i_exotiny._0369_[5] ),
    .A2(net1193));
 sg13g2_a21oi_1 _06727_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01408_),
    .A2(net1193),
    .Y(_02759_),
    .B1(_02758_));
 sg13g2_a221oi_1 _06728_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net8),
    .C1(_02759_),
    .B1(_02747_),
    .A1(net3795),
    .Y(_02760_),
    .A2(net1182));
 sg13g2_a221oi_1 _06729_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01506_),
    .C1(_02757_),
    .B1(_02760_),
    .A1(_01366_),
    .Y(_00665_),
    .A2(net1068));
 sg13g2_nand2_1 _06730_ (.Y(_02761_),
    .A(net3751),
    .B(net1183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06731_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01409_),
    .A2(net1192),
    .Y(_02762_),
    .B1(net1169));
 sg13g2_o21ai_1 _06732_ (.B1(_02762_),
    .VDD(VPWR),
    .Y(_02763_),
    .VSS(VGND),
    .A1(\i_exotiny._0369_[6] ),
    .A2(net1192));
 sg13g2_a21oi_1 _06733_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02761_),
    .A2(_02763_),
    .Y(_02764_),
    .B1(net1130));
 sg13g2_a21oi_1 _06734_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1980),
    .A2(net1137),
    .Y(_02765_),
    .B1(_02764_));
 sg13g2_nor2_1 _06735_ (.A(net3730),
    .B(net1101),
    .Y(_02766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06736_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1101),
    .A2(_02765_),
    .Y(_00666_),
    .B1(_02766_));
 sg13g2_nand2_1 _06737_ (.Y(_02767_),
    .A(net3714),
    .B(net1183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06738_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01410_),
    .A2(net1190),
    .Y(_02768_),
    .B1(net1169));
 sg13g2_o21ai_1 _06739_ (.B1(_02768_),
    .VDD(VPWR),
    .Y(_02769_),
    .VSS(VGND),
    .A1(\i_exotiny._0369_[7] ),
    .A2(net1192));
 sg13g2_a21oi_1 _06740_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02767_),
    .A2(_02769_),
    .Y(_02770_),
    .B1(net1130));
 sg13g2_a21oi_1 _06741_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2331),
    .A2(net1130),
    .Y(_02771_),
    .B1(_02770_));
 sg13g2_nor2_1 _06742_ (.A(net3611),
    .B(net1096),
    .Y(_02772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06743_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1101),
    .A2(_02771_),
    .Y(_00667_),
    .B1(_02772_));
 sg13g2_nand2_1 _06744_ (.Y(_02773_),
    .A(net3708),
    .B(net1183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06745_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01411_),
    .A2(net1190),
    .Y(_02774_),
    .B1(net1169));
 sg13g2_o21ai_1 _06746_ (.B1(_02774_),
    .VDD(VPWR),
    .Y(_02775_),
    .VSS(VGND),
    .A1(net3778),
    .A2(net1190));
 sg13g2_a21oi_1 _06747_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02773_),
    .A2(_02775_),
    .Y(_02776_),
    .B1(net1135));
 sg13g2_a21oi_1 _06748_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2042),
    .A2(net1130),
    .Y(_02777_),
    .B1(_02776_));
 sg13g2_nor2_1 _06749_ (.A(net3808),
    .B(net1100),
    .Y(_02778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06750_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1100),
    .A2(_02777_),
    .Y(_00668_),
    .B1(_02778_));
 sg13g2_o21ai_1 _06751_ (.B1(net1171),
    .VDD(VPWR),
    .Y(_02779_),
    .VSS(VGND),
    .A1(net1933),
    .A2(net1185));
 sg13g2_a21oi_1 _06752_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01406_),
    .A2(_01451_),
    .Y(_02780_),
    .B1(_02779_));
 sg13g2_a221oi_1 _06753_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net2106),
    .C1(_02780_),
    .B1(net3821),
    .A1(net3791),
    .Y(_02781_),
    .A2(net1182));
 sg13g2_a22oi_1 _06754_ (.Y(_02782_),
    .B1(_02719_),
    .B2(net3559),
    .A2(net1068),
    .A1(net3142),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06755_ (.B1(_02782_),
    .VDD(VPWR),
    .Y(_00669_),
    .VSS(VGND),
    .A1(net1137),
    .A2(_02781_));
 sg13g2_o21ai_1 _06756_ (.B1(net1171),
    .VDD(VPWR),
    .Y(_02783_),
    .VSS(VGND),
    .A1(net3443),
    .A2(net1191));
 sg13g2_a21oi_1 _06757_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01412_),
    .A2(net1191),
    .Y(_02784_),
    .B1(_02783_));
 sg13g2_a221oi_1 _06758_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net3656),
    .C1(_02784_),
    .B1(net3821),
    .A1(net3835),
    .Y(_02785_),
    .A2(net1182));
 sg13g2_or2_1 _06759_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_02786_),
    .B(net1102),
    .A(net1980));
 sg13g2_o21ai_1 _06760_ (.B1(_02786_),
    .VDD(VPWR),
    .Y(_02787_),
    .VSS(VGND),
    .A1(net3622),
    .A2(_02720_));
 sg13g2_a21oi_1 _06761_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01506_),
    .A2(_02785_),
    .Y(_00670_),
    .B1(_02787_));
 sg13g2_nand2_1 _06762_ (.Y(_02788_),
    .A(net1870),
    .B(net1183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06763_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01413_),
    .A2(net1190),
    .Y(_02789_),
    .B1(net1169));
 sg13g2_o21ai_1 _06764_ (.B1(_02789_),
    .VDD(VPWR),
    .Y(_02790_),
    .VSS(VGND),
    .A1(net3641),
    .A2(net1190));
 sg13g2_a21oi_1 _06765_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02788_),
    .A2(_02790_),
    .Y(_02791_),
    .B1(net1135));
 sg13g2_a21oi_1 _06766_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3801),
    .A2(net1135),
    .Y(_02792_),
    .B1(_02791_));
 sg13g2_nor2_1 _06767_ (.A(net2331),
    .B(net1100),
    .Y(_02793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06768_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1100),
    .A2(_02792_),
    .Y(_00671_),
    .B1(_02793_));
 sg13g2_nand2_1 _06769_ (.Y(_02794_),
    .A(net1875),
    .B(net1183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06770_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01414_),
    .A2(net1190),
    .Y(_02795_),
    .B1(net1169));
 sg13g2_o21ai_1 _06771_ (.B1(_02795_),
    .VDD(VPWR),
    .Y(_02796_),
    .VSS(VGND),
    .A1(net3759),
    .A2(net1190));
 sg13g2_a21oi_1 _06772_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02794_),
    .A2(_02796_),
    .Y(_02797_),
    .B1(net1135));
 sg13g2_a21oi_1 _06773_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2063),
    .A2(net1135),
    .Y(_02798_),
    .B1(_02797_));
 sg13g2_nor2_1 _06774_ (.A(net2042),
    .B(net1100),
    .Y(_02799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06775_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1100),
    .A2(_02798_),
    .Y(_00672_),
    .B1(_02799_));
 sg13g2_nand2_1 _06776_ (.Y(_02800_),
    .A(net1873),
    .B(net1183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06777_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01415_),
    .A2(net1192),
    .Y(_02801_),
    .B1(net1169));
 sg13g2_o21ai_1 _06778_ (.B1(_02801_),
    .VDD(VPWR),
    .Y(_02802_),
    .VSS(VGND),
    .A1(net3749),
    .A2(net1190));
 sg13g2_a21oi_1 _06779_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02800_),
    .A2(_02802_),
    .Y(_02803_),
    .B1(net1135));
 sg13g2_a21oi_1 _06780_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net2012),
    .A2(net1131),
    .Y(_02804_),
    .B1(_02803_));
 sg13g2_nor2_1 _06781_ (.A(net3559),
    .B(net1096),
    .Y(_02805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06782_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1096),
    .A2(_02804_),
    .Y(_00673_),
    .B1(_02805_));
 sg13g2_nor2_1 _06783_ (.A(net3643),
    .B(net1191),
    .Y(_02806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06784_ (.B1(net1171),
    .VDD(VPWR),
    .Y(_02807_),
    .VSS(VGND),
    .A1(net1945),
    .A2(_01451_));
 sg13g2_nor3_1 _06785_ (.A(net1132),
    .B(_02806_),
    .C(_02807_),
    .Y(_02808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06786_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3630),
    .A2(net1133),
    .Y(_02809_),
    .B1(_02808_));
 sg13g2_nor2_1 _06787_ (.A(net3622),
    .B(net1098),
    .Y(_02810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06788_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1098),
    .A2(_02809_),
    .Y(_00674_),
    .B1(_02810_));
 sg13g2_nor2_1 _06789_ (.A(net3596),
    .B(net1188),
    .Y(_02811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06790_ (.B1(net1171),
    .VDD(VPWR),
    .Y(_02812_),
    .VSS(VGND),
    .A1(net2432),
    .A2(net1185));
 sg13g2_nor3_1 _06791_ (.A(net1133),
    .B(_02811_),
    .C(_02812_),
    .Y(_02813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06792_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3711),
    .A2(net1133),
    .Y(_02814_),
    .B1(_02813_));
 sg13g2_nor2_1 _06793_ (.A(net3801),
    .B(net1098),
    .Y(_02815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06794_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1098),
    .A2(_02814_),
    .Y(_00675_),
    .B1(_02815_));
 sg13g2_nand2_1 _06795_ (.Y(_02816_),
    .A(net3733),
    .B(_02745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06796_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01416_),
    .A2(net1191),
    .Y(_02817_),
    .B1(_01517_));
 sg13g2_o21ai_1 _06797_ (.B1(_02817_),
    .VDD(VPWR),
    .Y(_02818_),
    .VSS(VGND),
    .A1(\i_exotiny._0369_[16] ),
    .A2(net1191));
 sg13g2_a21oi_1 _06798_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02816_),
    .A2(_02818_),
    .Y(_02819_),
    .B1(net1130));
 sg13g2_a21oi_1 _06799_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3717),
    .A2(net1130),
    .Y(_02820_),
    .B1(net3734));
 sg13g2_nor2_1 _06800_ (.A(net2063),
    .B(net1099),
    .Y(_02821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06801_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1099),
    .A2(_02820_),
    .Y(_00676_),
    .B1(_02821_));
 sg13g2_nand2_1 _06802_ (.Y(_02822_),
    .A(\i_exotiny.i_wb_regs.spi_size_o[1] ),
    .B(_02745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06803_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01417_),
    .A2(net1191),
    .Y(_02823_),
    .B1(_01517_));
 sg13g2_o21ai_1 _06804_ (.B1(_02823_),
    .VDD(VPWR),
    .Y(_02824_),
    .VSS(VGND),
    .A1(net3675),
    .A2(net1191));
 sg13g2_a21oi_1 _06805_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02822_),
    .A2(_02824_),
    .Y(_02825_),
    .B1(net1130));
 sg13g2_a21oi_1 _06806_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3697),
    .A2(net1130),
    .Y(_02826_),
    .B1(_02825_));
 sg13g2_nor2_1 _06807_ (.A(net2012),
    .B(net1096),
    .Y(_02827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06808_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1096),
    .A2(net3698),
    .Y(_00677_),
    .B1(_02827_));
 sg13g2_nor2_1 _06809_ (.A(\i_exotiny._0369_[18] ),
    .B(net1188),
    .Y(_02828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06810_ (.B1(net1171),
    .VDD(VPWR),
    .Y(_02829_),
    .VSS(VGND),
    .A1(net1937),
    .A2(net1185));
 sg13g2_nor3_1 _06811_ (.A(net1132),
    .B(_02828_),
    .C(_02829_),
    .Y(_02830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06812_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3563),
    .A2(net1132),
    .Y(_02831_),
    .B1(_02830_));
 sg13g2_nor2_1 _06813_ (.A(net3630),
    .B(net1097),
    .Y(_02832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06814_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1097),
    .A2(_02831_),
    .Y(_00678_),
    .B1(_02832_));
 sg13g2_nor2_1 _06815_ (.A(net3505),
    .B(net1189),
    .Y(_02833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06816_ (.B1(net1170),
    .VDD(VPWR),
    .Y(_02834_),
    .VSS(VGND),
    .A1(net3655),
    .A2(net1185));
 sg13g2_nor3_1 _06817_ (.A(net1132),
    .B(_02833_),
    .C(_02834_),
    .Y(_02835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06818_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3680),
    .A2(net1133),
    .Y(_02836_),
    .B1(_02835_));
 sg13g2_nor2_1 _06819_ (.A(net3711),
    .B(net1097),
    .Y(_02837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06820_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1097),
    .A2(_02836_),
    .Y(_00679_),
    .B1(_02837_));
 sg13g2_nor2_1 _06821_ (.A(\i_exotiny._0369_[20] ),
    .B(net1188),
    .Y(_02838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06822_ (.B1(net1170),
    .VDD(VPWR),
    .Y(_02839_),
    .VSS(VGND),
    .A1(net3644),
    .A2(net1185));
 sg13g2_nor3_1 _06823_ (.A(net1132),
    .B(_02838_),
    .C(_02839_),
    .Y(_02840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06824_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3501),
    .A2(net1134),
    .Y(_02841_),
    .B1(_02840_));
 sg13g2_nor2_1 _06825_ (.A(net3717),
    .B(net1099),
    .Y(_02842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06826_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1099),
    .A2(_02841_),
    .Y(_00680_),
    .B1(_02842_));
 sg13g2_nor2_1 _06827_ (.A(net2125),
    .B(net1188),
    .Y(_02843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06828_ (.B1(net1170),
    .VDD(VPWR),
    .Y(_02844_),
    .VSS(VGND),
    .A1(net3600),
    .A2(net1185));
 sg13g2_nor3_1 _06829_ (.A(net1132),
    .B(_02843_),
    .C(_02844_),
    .Y(_02845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06830_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3572),
    .A2(net1131),
    .Y(_02846_),
    .B1(_02845_));
 sg13g2_nor2_1 _06831_ (.A(net3697),
    .B(net1096),
    .Y(_02847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06832_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1096),
    .A2(_02846_),
    .Y(_00681_),
    .B1(_02847_));
 sg13g2_nor2_1 _06833_ (.A(net3307),
    .B(net1188),
    .Y(_02848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06834_ (.B1(net1170),
    .VDD(VPWR),
    .Y(_02849_),
    .VSS(VGND),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[22] ),
    .A2(net1185));
 sg13g2_nor3_1 _06835_ (.A(net1129),
    .B(_02848_),
    .C(_02849_),
    .Y(_02850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06836_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1616_[2] ),
    .A2(net1132),
    .Y(_02851_),
    .B1(_02850_));
 sg13g2_nor2_1 _06837_ (.A(net3563),
    .B(net1097),
    .Y(_02852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06838_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1097),
    .A2(_02851_),
    .Y(_00682_),
    .B1(_02852_));
 sg13g2_nor2_1 _06839_ (.A(net2061),
    .B(net1188),
    .Y(_02853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06840_ (.B1(net1170),
    .VDD(VPWR),
    .Y(_02854_),
    .VSS(VGND),
    .A1(net3638),
    .A2(net1185));
 sg13g2_nor3_1 _06841_ (.A(net1128),
    .B(_02853_),
    .C(_02854_),
    .Y(_02855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06842_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3620),
    .A2(net1132),
    .Y(_02856_),
    .B1(_02855_));
 sg13g2_nor2_1 _06843_ (.A(net3680),
    .B(net1097),
    .Y(_02857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06844_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1097),
    .A2(_02856_),
    .Y(_00683_),
    .B1(_02857_));
 sg13g2_nor2_1 _06845_ (.A(\i_exotiny._0369_[24] ),
    .B(net1188),
    .Y(_02858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06846_ (.B1(net1170),
    .VDD(VPWR),
    .Y(_02859_),
    .VSS(VGND),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[24] ),
    .A2(net1186));
 sg13g2_nor3_1 _06847_ (.A(net1129),
    .B(_02858_),
    .C(_02859_),
    .Y(_02860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06848_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1619_[0] ),
    .A2(net1134),
    .Y(_02861_),
    .B1(_02860_));
 sg13g2_nor2_1 _06849_ (.A(net3501),
    .B(net1099),
    .Y(_02862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1094),
    .A2(_02861_),
    .Y(_00684_),
    .B1(_02862_));
 sg13g2_nor2_1 _06851_ (.A(\i_exotiny._0369_[25] ),
    .B(net1189),
    .Y(_02863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06852_ (.B1(net1170),
    .VDD(VPWR),
    .Y(_02864_),
    .VSS(VGND),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[25] ),
    .A2(net1186));
 sg13g2_nor3_1 _06853_ (.A(net1129),
    .B(_02863_),
    .C(_02864_),
    .Y(_02865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06854_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1619_[1] ),
    .A2(net1131),
    .Y(_02866_),
    .B1(_02865_));
 sg13g2_nor2_1 _06855_ (.A(net3572),
    .B(net1096),
    .Y(_02867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06856_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1094),
    .A2(_02866_),
    .Y(_00685_),
    .B1(_02867_));
 sg13g2_nor2_1 _06857_ (.A(net1872),
    .B(net1189),
    .Y(_02868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06858_ (.B1(net1171),
    .VDD(VPWR),
    .Y(_02869_),
    .VSS(VGND),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[26] ),
    .A2(net1186));
 sg13g2_nor3_1 _06859_ (.A(net1129),
    .B(_02868_),
    .C(_02869_),
    .Y(_02870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06860_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1619_[2] ),
    .A2(net1134),
    .Y(_02871_),
    .B1(_02870_));
 sg13g2_nor2_1 _06861_ (.A(net3614),
    .B(net1095),
    .Y(_02872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06862_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1095),
    .A2(_02871_),
    .Y(_00686_),
    .B1(_02872_));
 sg13g2_nor2_1 _06863_ (.A(net3584),
    .B(net1188),
    .Y(_02873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06864_ (.B1(net1170),
    .VDD(VPWR),
    .Y(_02874_),
    .VSS(VGND),
    .A1(net3616),
    .A2(net1186));
 sg13g2_nor3_1 _06865_ (.A(net1129),
    .B(_02873_),
    .C(_02874_),
    .Y(_02875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06866_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1619_[3] ),
    .A2(net1134),
    .Y(_02876_),
    .B1(_02875_));
 sg13g2_nor2_1 _06867_ (.A(net3620),
    .B(net1095),
    .Y(_02877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06868_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1095),
    .A2(_02876_),
    .Y(_00687_),
    .B1(_02877_));
 sg13g2_nor2_1 _06869_ (.A(\i_exotiny._0369_[28] ),
    .B(net1189),
    .Y(_02878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06870_ (.B1(net1172),
    .VDD(VPWR),
    .Y(_02879_),
    .VSS(VGND),
    .A1(net3623),
    .A2(net1186));
 sg13g2_nor3_1 _06871_ (.A(net1128),
    .B(_02878_),
    .C(_02879_),
    .Y(_02880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06872_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1618_[0] ),
    .A2(net1128),
    .Y(_02881_),
    .B1(_02880_));
 sg13g2_nor2_1 _06873_ (.A(net3668),
    .B(net1094),
    .Y(_02882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06874_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1094),
    .A2(_02881_),
    .Y(_00688_),
    .B1(_02882_));
 sg13g2_nor2_1 _06875_ (.A(net3601),
    .B(net1189),
    .Y(_02883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06876_ (.B1(net1172),
    .VDD(VPWR),
    .Y(_02884_),
    .VSS(VGND),
    .A1(net3646),
    .A2(net1186));
 sg13g2_nor3_1 _06877_ (.A(net1128),
    .B(_02883_),
    .C(_02884_),
    .Y(_02885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06878_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3422),
    .A2(net1131),
    .Y(_02886_),
    .B1(_02885_));
 sg13g2_nor2_1 _06879_ (.A(net3687),
    .B(net1094),
    .Y(_02887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06880_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1094),
    .A2(_02886_),
    .Y(_00689_),
    .B1(_02887_));
 sg13g2_nor2_1 _06881_ (.A(net3457),
    .B(net1189),
    .Y(_02888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06882_ (.B1(net1172),
    .VDD(VPWR),
    .Y(_02889_),
    .VSS(VGND),
    .A1(net3582),
    .A2(net1186));
 sg13g2_nor3_1 _06883_ (.A(net1128),
    .B(_02888_),
    .C(_02889_),
    .Y(_02890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06884_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1618_[2] ),
    .A2(net1128),
    .Y(_02891_),
    .B1(_02890_));
 sg13g2_nor2_1 _06885_ (.A(net3672),
    .B(net1094),
    .Y(_02892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06886_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1094),
    .A2(_02891_),
    .Y(_00690_),
    .B1(_02892_));
 sg13g2_nor2_1 _06887_ (.A(net3387),
    .B(net1189),
    .Y(_02893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06888_ (.B1(net1172),
    .VDD(VPWR),
    .Y(_02894_),
    .VSS(VGND),
    .A1(net3530),
    .A2(net1186));
 sg13g2_nor3_1 _06889_ (.A(net1128),
    .B(_02893_),
    .C(_02894_),
    .Y(_02895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06890_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1618_[3] ),
    .A2(net1128),
    .Y(_02896_),
    .B1(_02895_));
 sg13g2_nor2_1 _06891_ (.A(net3747),
    .B(net1095),
    .Y(_02897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06892_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1095),
    .A2(_02896_),
    .Y(_00691_),
    .B1(_02897_));
 sg13g2_a22oi_1 _06893_ (.Y(_02898_),
    .B1(_02719_),
    .B2(_02437_),
    .A2(net1068),
    .A1(net3811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _06894_ (.VDD(VPWR),
    .Y(_00692_),
    .A(_02898_),
    .VSS(VGND));
 sg13g2_nand2_1 _06895_ (.Y(_02899_),
    .A(net3422),
    .B(net1068),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _06896_ (.B1(_02899_),
    .VDD(VPWR),
    .Y(_00693_),
    .VSS(VGND),
    .A1(_02453_),
    .A2(_02720_));
 sg13g2_a22oi_1 _06897_ (.Y(_02900_),
    .B1(_02719_),
    .B2(_02462_),
    .A2(net1068),
    .A1(net3817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _06898_ (.VDD(VPWR),
    .Y(_00694_),
    .A(_02900_),
    .VSS(VGND));
 sg13g2_a22oi_1 _06899_ (.Y(_02901_),
    .B1(_02719_),
    .B2(_02471_),
    .A2(net1068),
    .A1(net3816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _06900_ (.VDD(VPWR),
    .Y(_00695_),
    .A(_02901_),
    .VSS(VGND));
 sg13g2_nand2b_1 _06901_ (.Y(_02902_),
    .B(net1970),
    .A_N(net3766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _06902_ (.A(net3658),
    .B(net2298),
    .C(net3681),
    .D(_02902_),
    .Y(_02903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06903_ (.Y(_02904_),
    .A(net3241),
    .B(net3466),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _06904_ (.A(net2570),
    .B(net1883),
    .C(_01389_),
    .D(_02904_),
    .Y(_02905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06905_ (.A2(_02905_),
    .A1(_02903_),
    .B1(net1227),
    .X(_02906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06906_ (.Y(_02907_),
    .A(net2570),
    .B(net1263),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _06907_ (.B(net2570),
    .C(net1263),
    .A(net3241),
    .Y(_02908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06908_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01368_),
    .A2(_02908_),
    .Y(_00696_),
    .B1(_02906_));
 sg13g2_nand2_1 _06909_ (.Y(_02909_),
    .A(\i_exotiny._1586_ ),
    .B(\i_exotiny.i_rstctl.cnt[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _06910_ (.B(\i_exotiny.i_rstctl.cnt[1] ),
    .C(\i_exotiny.i_rstctl.cnt[5] ),
    .A(net1883),
    .Y(_02910_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\i_exotiny.i_rstctl.cnt[4] ));
 sg13g2_nor4_1 _06911_ (.A(net2298),
    .B(net1970),
    .C(_02909_),
    .D(_02910_),
    .Y(_02911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06912_ (.A2(net3466),
    .A1(\i_exotiny.core_res_en_n ),
    .B1(_02911_),
    .X(_02912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _06913_ (.B(_01389_),
    .C(net3682),
    .A(net1883),
    .Y(_02913_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02912_));
 sg13g2_a21o_1 _06914_ (.A2(net3683),
    .A1(net2570),
    .B1(_02906_),
    .X(_00697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _06915_ (.Y(_02914_),
    .A(net2570),
    .B(_02912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _06916_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.core_res_en_n ),
    .A2(_02907_),
    .Y(_02915_),
    .B1(net1227));
 sg13g2_nand2_1 _06917_ (.Y(_00698_),
    .A(net2571),
    .B(_02915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06918_ (.A(_02485_),
    .B(_02532_),
    .Y(_02916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _06919_ (.A2(_02916_),
    .A1(net1138),
    .B1(net1165),
    .X(_02917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06920_ (.A0(\i_exotiny._0029_[0] ),
    .A1(net2635),
    .S(net926),
    .X(_00699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06921_ (.A0(\i_exotiny._0029_[1] ),
    .A1(net2524),
    .S(net924),
    .X(_00700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06922_ (.A0(\i_exotiny._0029_[2] ),
    .A1(net2408),
    .S(net926),
    .X(_00701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06923_ (.A0(net2720),
    .A1(net2721),
    .S(net927),
    .X(_00702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06924_ (.A0(net2635),
    .A1(net2688),
    .S(net926),
    .X(_00703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06925_ (.A0(net2524),
    .A1(net2856),
    .S(net924),
    .X(_00704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06926_ (.A0(net2408),
    .A1(net2783),
    .S(net925),
    .X(_00705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06927_ (.A0(net2721),
    .A1(net2848),
    .S(net927),
    .X(_00706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06928_ (.A0(net2688),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[12] ),
    .S(net926),
    .X(_00707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06929_ (.A0(net2856),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[13] ),
    .S(net924),
    .X(_00708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06930_ (.A0(net2783),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[14] ),
    .S(net925),
    .X(_00709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06931_ (.A0(net2848),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[15] ),
    .S(net927),
    .X(_00710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06932_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[12] ),
    .A1(net3380),
    .S(net926),
    .X(_00711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06933_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[13] ),
    .A1(net2265),
    .S(net924),
    .X(_00712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06934_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[14] ),
    .A1(net3299),
    .S(net925),
    .X(_00713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06935_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[15] ),
    .A1(net3041),
    .S(net927),
    .X(_00714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06936_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[16] ),
    .A1(net3032),
    .S(net926),
    .X(_00715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06937_ (.A0(net2265),
    .A1(net2503),
    .S(net924),
    .X(_00716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06938_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[18] ),
    .A1(net2278),
    .S(net925),
    .X(_00717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06939_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[19] ),
    .A1(net2315),
    .S(net927),
    .X(_00718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06940_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[20] ),
    .A1(net2192),
    .S(net928),
    .X(_00719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06941_ (.A0(net2503),
    .A1(net2747),
    .S(net924),
    .X(_00720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06942_ (.A0(net2278),
    .A1(net3056),
    .S(net925),
    .X(_00721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06943_ (.A0(net2315),
    .A1(net2488),
    .S(net927),
    .X(_00722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06944_ (.A0(net2192),
    .A1(net2734),
    .S(net926),
    .X(_00723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06945_ (.A0(net2747),
    .A1(net2897),
    .S(net924),
    .X(_00724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06946_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[26] ),
    .A1(net2927),
    .S(net925),
    .X(_00725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06947_ (.A0(net2488),
    .A1(net2575),
    .S(net927),
    .X(_00726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06948_ (.A0(net2985),
    .A1(net887),
    .S(_02916_),
    .X(_02918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06949_ (.A0(net2734),
    .A1(_02918_),
    .S(net926),
    .X(_00727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06950_ (.A0(net3187),
    .A1(net882),
    .S(_02916_),
    .X(_02919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06951_ (.A0(net2897),
    .A1(_02919_),
    .S(net924),
    .X(_00728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06952_ (.A0(net3043),
    .A1(net877),
    .S(_02916_),
    .X(_02920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06953_ (.A0(net2927),
    .A1(_02920_),
    .S(net925),
    .X(_00729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06954_ (.A0(net2720),
    .A1(net873),
    .S(_02916_),
    .X(_02921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06955_ (.A0(net2575),
    .A1(_02921_),
    .S(net927),
    .X(_00730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06956_ (.A(_02492_),
    .B(_02518_),
    .Y(_02922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _06957_ (.A2(_02922_),
    .A1(net1140),
    .B1(net1167),
    .X(_02923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06958_ (.A0(net2450),
    .A1(net3436),
    .S(net1021),
    .X(_00731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06959_ (.A0(\i_exotiny._0034_[1] ),
    .A1(net2677),
    .S(net1018),
    .X(_00732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06960_ (.A0(\i_exotiny._0034_[2] ),
    .A1(net2243),
    .S(net1022),
    .X(_00733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06961_ (.A0(net2805),
    .A1(net3247),
    .S(net1019),
    .X(_00734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06962_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[4] ),
    .A1(net3309),
    .S(net1021),
    .X(_00735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06963_ (.A0(net2677),
    .A1(net2944),
    .S(net1018),
    .X(_00736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06964_ (.A0(net2243),
    .A1(net3372),
    .S(net1022),
    .X(_00737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06965_ (.A0(net3247),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[11] ),
    .S(net1019),
    .X(_00738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06966_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[8] ),
    .A1(net3099),
    .S(net1021),
    .X(_00739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06967_ (.A0(net2944),
    .A1(net2988),
    .S(net1018),
    .X(_00740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06968_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[10] ),
    .A1(net3216),
    .S(net1020),
    .X(_00741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06969_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[11] ),
    .A1(net3288),
    .S(net1020),
    .X(_00742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06970_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[12] ),
    .A1(net2722),
    .S(net1021),
    .X(_00743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06971_ (.A0(net2988),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[17] ),
    .S(net1018),
    .X(_00744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06972_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[14] ),
    .A1(net2329),
    .S(net1020),
    .X(_00745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06973_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[15] ),
    .A1(net2280),
    .S(net1020),
    .X(_00746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06974_ (.A0(net2722),
    .A1(net2908),
    .S(net1021),
    .X(_00747_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06975_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[17] ),
    .A1(net1994),
    .S(net1018),
    .X(_00748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06976_ (.A0(net2329),
    .A1(net2819),
    .S(net1022),
    .X(_00749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06977_ (.A0(net2280),
    .A1(net2945),
    .S(net1020),
    .X(_00750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06978_ (.A0(net2908),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[24] ),
    .S(net1021),
    .X(_00751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06979_ (.A0(net1994),
    .A1(net2656),
    .S(net1018),
    .X(_00752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06980_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[22] ),
    .A1(net2770),
    .S(net1020),
    .X(_00753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06981_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[23] ),
    .A1(net2925),
    .S(net1019),
    .X(_00754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06982_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[24] ),
    .A1(net2355),
    .S(net1021),
    .X(_00755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06983_ (.A0(net2656),
    .A1(net2742),
    .S(net1018),
    .X(_00756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06984_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[26] ),
    .A1(net2160),
    .S(net1020),
    .X(_00757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06985_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[27] ),
    .A1(net2178),
    .S(net1019),
    .X(_00758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06986_ (.A0(net2450),
    .A1(net889),
    .S(_02922_),
    .X(_02924_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06987_ (.A0(net2355),
    .A1(_02924_),
    .S(net1021),
    .X(_00759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06988_ (.A0(net3104),
    .A1(net883),
    .S(_02922_),
    .X(_02925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06989_ (.A0(net2742),
    .A1(_02925_),
    .S(net1018),
    .X(_00760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06990_ (.A0(net2803),
    .A1(net879),
    .S(_02922_),
    .X(_02926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06991_ (.A0(net2160),
    .A1(_02926_),
    .S(net1020),
    .X(_00761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06992_ (.A0(net2805),
    .A1(net875),
    .S(_02922_),
    .X(_02927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06993_ (.A0(net2178),
    .A1(_02927_),
    .S(net1019),
    .X(_00762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _06994_ (.A(_02517_),
    .B(_02532_),
    .Y(_02928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _06995_ (.A2(_02928_),
    .A1(net1141),
    .B1(net1165),
    .X(_02929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06996_ (.A0(\i_exotiny._0032_[0] ),
    .A1(net2059),
    .S(net922),
    .X(_00763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06997_ (.A0(net3202),
    .A1(net3497),
    .S(net920),
    .X(_00764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06998_ (.A0(\i_exotiny._0032_[2] ),
    .A1(net2627),
    .S(net919),
    .X(_00765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _06999_ (.A0(\i_exotiny._0032_[3] ),
    .A1(net2093),
    .S(net918),
    .X(_00766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07000_ (.A0(net2059),
    .A1(net2765),
    .S(net922),
    .X(_00767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07001_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[5] ),
    .A1(net2089),
    .S(net920),
    .X(_00768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07002_ (.A0(net2627),
    .A1(net3178),
    .S(net919),
    .X(_00769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07003_ (.A0(net2093),
    .A1(net2972),
    .S(net918),
    .X(_00770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07004_ (.A0(net2765),
    .A1(net2872),
    .S(net922),
    .X(_00771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07005_ (.A0(net2089),
    .A1(net3028),
    .S(net920),
    .X(_00772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07006_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[10] ),
    .A1(net3034),
    .S(net921),
    .X(_00773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07007_ (.A0(net2972),
    .A1(net3130),
    .S(net918),
    .X(_00774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07008_ (.A0(net2872),
    .A1(net2645),
    .S(net922),
    .X(_00775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07009_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[13] ),
    .A1(net2075),
    .S(net921),
    .X(_00776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07010_ (.A0(net3034),
    .A1(net3093),
    .S(net921),
    .X(_00777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07011_ (.A0(net3130),
    .A1(net2912),
    .S(net918),
    .X(_00778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07012_ (.A0(net2645),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[20] ),
    .S(net922),
    .X(_00779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07013_ (.A0(net2075),
    .A1(net2746),
    .S(net921),
    .X(_00780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07014_ (.A0(net3093),
    .A1(net3287),
    .S(net920),
    .X(_00781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07015_ (.A0(net2912),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[23] ),
    .S(net918),
    .X(_00782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07016_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[20] ),
    .A1(net3395),
    .S(net922),
    .X(_00783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07017_ (.A0(net2746),
    .A1(net2994),
    .S(net921),
    .X(_00784_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07018_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[22] ),
    .A1(net2111),
    .S(net920),
    .X(_00785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07019_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[23] ),
    .A1(net3183),
    .S(net918),
    .X(_00786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07020_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[24] ),
    .A1(net2083),
    .S(net922),
    .X(_00787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07021_ (.A0(net2994),
    .A1(net3175),
    .S(net920),
    .X(_00788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07022_ (.A0(net2111),
    .A1(net3077),
    .S(net920),
    .X(_00789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07023_ (.A0(net3183),
    .A1(net3301),
    .S(net918),
    .X(_00790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07024_ (.A0(net3320),
    .A1(net887),
    .S(_02928_),
    .X(_02930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07025_ (.A0(net2083),
    .A1(_02930_),
    .S(net918),
    .X(_00791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07026_ (.A0(net3202),
    .A1(net884),
    .S(_02928_),
    .X(_02931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07027_ (.A0(net3175),
    .A1(_02931_),
    .S(net920),
    .X(_00792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07028_ (.A0(\i_exotiny._0032_[2] ),
    .A1(net877),
    .S(_02928_),
    .X(_02932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07029_ (.A0(net3077),
    .A1(_02932_),
    .S(net919),
    .X(_00793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07030_ (.A0(net3452),
    .A1(net875),
    .S(_02928_),
    .X(_02933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07031_ (.A0(net3301),
    .A1(_02933_),
    .S(net919),
    .X(_00794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07032_ (.A(_02420_),
    .B(_02564_),
    .Y(_02934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _07033_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net1166),
    .Y(_02935_),
    .A2(_02934_),
    .A1(net1139));
 sg13g2_mux2_1 _07034_ (.A0(net2410),
    .A1(\i_exotiny._0017_[0] ),
    .S(net1013),
    .X(_00795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07035_ (.A0(net3593),
    .A1(net3129),
    .S(net1014),
    .X(_00796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07036_ (.A0(net3356),
    .A1(net2866),
    .S(net1017),
    .X(_00797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07037_ (.A0(net3109),
    .A1(net3065),
    .S(net1014),
    .X(_00798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07038_ (.A0(net2548),
    .A1(net2410),
    .S(net1013),
    .X(_00799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07039_ (.A0(net2293),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[5] ),
    .S(net1015),
    .X(_00800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07040_ (.A0(net2920),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[6] ),
    .S(net1017),
    .X(_00801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07041_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[11] ),
    .A1(net3109),
    .S(net1013),
    .X(_00802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07042_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[12] ),
    .A1(net2548),
    .S(net1013),
    .X(_00803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07043_ (.A0(net1828),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[9] ),
    .S(net1015),
    .X(_00804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07044_ (.A0(net3194),
    .A1(net2920),
    .S(net1017),
    .X(_00805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07045_ (.A0(net3199),
    .A1(net3449),
    .S(net1016),
    .X(_00806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07046_ (.A0(net2393),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[12] ),
    .S(net1013),
    .X(_00807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07047_ (.A0(net2222),
    .A1(net1828),
    .S(net1015),
    .X(_00808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07048_ (.A0(net3045),
    .A1(net3194),
    .S(net1017),
    .X(_00809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07049_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[19] ),
    .A1(net3199),
    .S(net1016),
    .X(_00810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07050_ (.A0(net3255),
    .A1(net2393),
    .S(net1014),
    .X(_00811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07051_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[21] ),
    .A1(net2222),
    .S(net1015),
    .X(_00812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07052_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[22] ),
    .A1(net3045),
    .S(net1017),
    .X(_00813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07053_ (.A0(net3425),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[19] ),
    .S(net1015),
    .X(_00814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07054_ (.A0(net2830),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[20] ),
    .S(net1013),
    .X(_00815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07055_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[25] ),
    .A1(net2573),
    .S(net1015),
    .X(_00816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07056_ (.A0(net3275),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[22] ),
    .S(net1017),
    .X(_00817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07057_ (.A0(net2555),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[23] ),
    .S(net1016),
    .X(_00818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07058_ (.A0(net3304),
    .A1(net2830),
    .S(net1013),
    .X(_00819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07059_ (.A0(net2806),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[25] ),
    .S(net1015),
    .X(_00820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07060_ (.A0(net2313),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[26] ),
    .S(net1017),
    .X(_00821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07061_ (.A0(net3047),
    .A1(net2555),
    .S(net1015),
    .X(_00822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07062_ (.A0(\i_exotiny._0017_[0] ),
    .A1(net888),
    .S(_02934_),
    .X(_02936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07063_ (.A0(_02936_),
    .A1(net3304),
    .S(net1013),
    .X(_00823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07064_ (.A0(net3129),
    .A1(net883),
    .S(_02934_),
    .X(_02937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07065_ (.A0(_02937_),
    .A1(net2806),
    .S(net1014),
    .X(_00824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07066_ (.A0(net2866),
    .A1(net878),
    .S(_02934_),
    .X(_02938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07067_ (.A0(_02938_),
    .A1(net2313),
    .S(net1017),
    .X(_00825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07068_ (.A0(net3065),
    .A1(net874),
    .S(_02934_),
    .X(_02939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07069_ (.A0(_02939_),
    .A1(net3047),
    .S(net1014),
    .X(_00826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07070_ (.A(_02420_),
    .B(_02517_),
    .Y(_02940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07071_ (.A2(_02940_),
    .A1(net1142),
    .B1(net1163),
    .X(_02941_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07072_ (.A0(net3063),
    .A1(net3000),
    .S(net914),
    .X(_00827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07073_ (.A0(\i_exotiny._0015_[1] ),
    .A1(net3368),
    .S(net916),
    .X(_00828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07074_ (.A0(net3080),
    .A1(net3073),
    .S(net916),
    .X(_00829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07075_ (.A0(\i_exotiny._0015_[3] ),
    .A1(net2359),
    .S(net916),
    .X(_00830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07076_ (.A0(net3000),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[8] ),
    .S(net914),
    .X(_00831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07077_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[5] ),
    .A1(net3039),
    .S(net916),
    .X(_00832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07078_ (.A0(net3073),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[10] ),
    .S(net916),
    .X(_00833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07079_ (.A0(net2359),
    .A1(net2644),
    .S(net915),
    .X(_00834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07080_ (.A0(net3335),
    .A1(net3076),
    .S(net913),
    .X(_00835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07081_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[9] ),
    .A1(net2144),
    .S(net913),
    .X(_00836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07082_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[10] ),
    .A1(net3364),
    .S(net916),
    .X(_00837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07083_ (.A0(net2644),
    .A1(net3404),
    .S(net915),
    .X(_00838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07084_ (.A0(net3076),
    .A1(net2967),
    .S(net913),
    .X(_00839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07085_ (.A0(net2144),
    .A1(net3197),
    .S(net913),
    .X(_00840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07086_ (.A0(net3364),
    .A1(net3367),
    .S(net917),
    .X(_00841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07087_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[15] ),
    .A1(net3330),
    .S(net915),
    .X(_00842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07088_ (.A0(net2967),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[20] ),
    .S(net913),
    .X(_00843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07089_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[17] ),
    .A1(net2158),
    .S(net915),
    .X(_00844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07090_ (.A0(net3367),
    .A1(net3440),
    .S(net917),
    .X(_00845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07091_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[19] ),
    .A1(net2117),
    .S(net914),
    .X(_00846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07092_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[20] ),
    .A1(net3413),
    .S(net913),
    .X(_00847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07093_ (.A0(net2158),
    .A1(net2512),
    .S(net915),
    .X(_00848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07094_ (.A0(net3440),
    .A1(net3464),
    .S(net916),
    .X(_00849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07095_ (.A0(net2117),
    .A1(net2289),
    .S(net914),
    .X(_00850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07096_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[24] ),
    .A1(net2694),
    .S(net914),
    .X(_00851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07097_ (.A0(net2512),
    .A1(net2936),
    .S(net913),
    .X(_00852_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07098_ (.A0(net3464),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[30] ),
    .S(net917),
    .X(_00853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07099_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[27] ),
    .A1(net2216),
    .S(net914),
    .X(_00854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07100_ (.A0(net3063),
    .A1(net886),
    .S(_02940_),
    .X(_02942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07101_ (.A0(net2694),
    .A1(_02942_),
    .S(net914),
    .X(_00855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07102_ (.A0(\i_exotiny._0015_[1] ),
    .A1(net881),
    .S(_02940_),
    .X(_02943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07103_ (.A0(net2936),
    .A1(_02943_),
    .S(net913),
    .X(_00856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07104_ (.A0(net3080),
    .A1(net876),
    .S(_02940_),
    .X(_02944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07105_ (.A0(net3507),
    .A1(_02944_),
    .S(net916),
    .X(_00857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07106_ (.A0(net3002),
    .A1(net872),
    .S(_02940_),
    .X(_02945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07107_ (.A0(net2216),
    .A1(_02945_),
    .S(net914),
    .X(_00858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07108_ (.A2(_02381_),
    .A1(net1111),
    .B1(net1227),
    .X(_02946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07109_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01379_),
    .A2(_01579_),
    .Y(_00859_),
    .B1(_02946_));
 sg13g2_and2_1 _07110_ (.A(net1288),
    .B(net1863),
    .X(_00860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07111_ (.A(net1288),
    .B(net1861),
    .X(_00861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07112_ (.A(net1288),
    .B(net1851),
    .X(_00862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07113_ (.A(net1286),
    .B(net1869),
    .X(_00863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07114_ (.A(net1288),
    .B(net1848),
    .X(_00864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07115_ (.A(net1289),
    .B(net1855),
    .X(_00865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07116_ (.A(net1289),
    .B(net1857),
    .X(_00866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07117_ (.A(net1288),
    .B(net1846),
    .X(_00867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07118_ (.A(net1288),
    .B(net1847),
    .X(_00868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07119_ (.A(net1288),
    .B(net1853),
    .X(_00869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07120_ (.A(net1288),
    .B(net1858),
    .X(_00870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07121_ (.A(net1290),
    .B(net1849),
    .X(_00871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07122_ (.A(net1289),
    .B(net1837),
    .X(_00872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07123_ (.A(net1290),
    .B(net1835),
    .X(_00873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07124_ (.A(net1290),
    .B(net1841),
    .X(_00874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07125_ (.A(net1287),
    .B(net1867),
    .X(_00875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07126_ (.A(net1290),
    .B(net1859),
    .X(_00876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07127_ (.A(net1287),
    .B(net1865),
    .X(_00877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07128_ (.A(net1287),
    .B(net1868),
    .X(_00878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07129_ (.A(net1287),
    .B(net1852),
    .X(_00879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07130_ (.A(net1289),
    .B(net1839),
    .X(_00880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07131_ (.A(net1287),
    .B(net1856),
    .X(_00881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07132_ (.A(net1287),
    .B(net1845),
    .X(_00882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07133_ (.A(net1286),
    .B(net1862),
    .X(_00883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07134_ (.A(net1287),
    .B(net1843),
    .X(_00884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07135_ (.A(net1286),
    .B(net1834),
    .X(_00885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07136_ (.A(net1286),
    .B(net1838),
    .X(_00886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07137_ (.A(net1286),
    .B(net1866),
    .X(_00887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07138_ (.A(net1286),
    .B(net1844),
    .X(_00888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07139_ (.A(net1286),
    .B(net1864),
    .X(_00889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07140_ (.A(net1286),
    .B(net1854),
    .X(_00890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07141_ (.A(_02419_),
    .B(_02532_),
    .Y(_02947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _07142_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net1159),
    .Y(_02948_),
    .A2(_02947_),
    .A1(net1142));
 sg13g2_mux2_1 _07143_ (.A0(net2174),
    .A1(\i_exotiny._0036_[0] ),
    .S(net1011),
    .X(_00891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07144_ (.A0(net2204),
    .A1(\i_exotiny._0036_[1] ),
    .S(net1012),
    .X(_00892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07145_ (.A0(net3281),
    .A1(net3397),
    .S(net1012),
    .X(_00893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07146_ (.A0(net2079),
    .A1(\i_exotiny._0036_[3] ),
    .S(net1012),
    .X(_00894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07147_ (.A0(net2652),
    .A1(net2174),
    .S(net1011),
    .X(_00895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07148_ (.A0(net2828),
    .A1(net2204),
    .S(net1012),
    .X(_00896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07149_ (.A0(net2787),
    .A1(net3281),
    .S(net1011),
    .X(_00897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07150_ (.A0(net2858),
    .A1(net2079),
    .S(net1012),
    .X(_00898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07151_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[12] ),
    .A1(net2652),
    .S(net1012),
    .X(_00899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07152_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[13] ),
    .A1(net2828),
    .S(net1009),
    .X(_00900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07153_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[14] ),
    .A1(net2787),
    .S(net1010),
    .X(_00901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07154_ (.A0(net3107),
    .A1(net2858),
    .S(net1009),
    .X(_00902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07155_ (.A0(net2323),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[12] ),
    .S(net1011),
    .X(_00903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07156_ (.A0(net2198),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[13] ),
    .S(net1008),
    .X(_00904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07157_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[18] ),
    .A1(net3214),
    .S(net1010),
    .X(_00905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07158_ (.A0(net3016),
    .A1(net3107),
    .S(net1008),
    .X(_00906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07159_ (.A0(net3167),
    .A1(net2323),
    .S(net1011),
    .X(_00907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07160_ (.A0(net2213),
    .A1(net2198),
    .S(net1008),
    .X(_00908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07161_ (.A0(net2052),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[18] ),
    .S(net1010),
    .X(_00909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07162_ (.A0(net2442),
    .A1(net3016),
    .S(net1008),
    .X(_00910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07163_ (.A0(net2711),
    .A1(net3167),
    .S(net1012),
    .X(_00911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07164_ (.A0(net3160),
    .A1(net2213),
    .S(net1008),
    .X(_00912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07165_ (.A0(net2608),
    .A1(net2052),
    .S(net1010),
    .X(_00913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07166_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[27] ),
    .A1(net2442),
    .S(net1009),
    .X(_00914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07167_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[28] ),
    .A1(net2711),
    .S(net1011),
    .X(_00915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07168_ (.A0(net2660),
    .A1(net3160),
    .S(net1008),
    .X(_00916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07169_ (.A0(net2861),
    .A1(net2608),
    .S(net1010),
    .X(_00917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07170_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[31] ),
    .A1(net2956),
    .S(net1008),
    .X(_00918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07171_ (.A0(\i_exotiny._0036_[0] ),
    .A1(net886),
    .S(_02947_),
    .X(_02949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07172_ (.A0(_02949_),
    .A1(net3533),
    .S(net1011),
    .X(_00919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07173_ (.A0(\i_exotiny._0036_[1] ),
    .A1(net881),
    .S(_02947_),
    .X(_02950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07174_ (.A0(_02950_),
    .A1(net2660),
    .S(net1008),
    .X(_00920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07175_ (.A0(net3397),
    .A1(net876),
    .S(_02947_),
    .X(_02951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07176_ (.A0(_02951_),
    .A1(net2861),
    .S(net1011),
    .X(_00921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07177_ (.A0(\i_exotiny._0036_[3] ),
    .A1(net872),
    .S(_02947_),
    .X(_02952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07178_ (.A0(_02952_),
    .A1(net3437),
    .S(net1009),
    .X(_00922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07179_ (.A(_02126_),
    .B(_02596_),
    .Y(_02953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07180_ (.Y(_02954_),
    .A(net1285),
    .B(_02953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07181_ (.A0(net3622),
    .A1(net3656),
    .S(_02954_),
    .X(_00923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07182_ (.Y(_02955_),
    .A(net2106),
    .B(net1285),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07183_ (.Y(_00924_),
    .B1(_02954_),
    .B2(net2107),
    .A2(_02953_),
    .A1(_01367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _07184_ (.A(net3762),
    .B(net1233),
    .C(\i_exotiny._0315_[4] ),
    .Y(_02956_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_02594_));
 sg13g2_o21ai_1 _07185_ (.B1(net1281),
    .VDD(VPWR),
    .Y(_02957_),
    .VSS(VGND),
    .A1(net3772),
    .A2(_02956_));
 sg13g2_a21oi_1 _07186_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01361_),
    .A2(_02956_),
    .Y(_00925_),
    .B1(net3773));
 sg13g2_o21ai_1 _07187_ (.B1(net1281),
    .VDD(VPWR),
    .Y(_02958_),
    .VSS(VGND),
    .A1(net3741),
    .A2(_02956_));
 sg13g2_a21oi_1 _07188_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01366_),
    .A2(_02956_),
    .Y(_00926_),
    .B1(net3742));
 sg13g2_o21ai_1 _07189_ (.B1(net1281),
    .VDD(VPWR),
    .Y(_02959_),
    .VSS(VGND),
    .A1(net3744),
    .A2(_02956_));
 sg13g2_a21oi_1 _07190_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01365_),
    .A2(_02956_),
    .Y(_00927_),
    .B1(net3745));
 sg13g2_nand2_1 _07191_ (.Y(_02960_),
    .A(net3606),
    .B(net1111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07192_ (.A0(net9),
    .A1(net3589),
    .S(net1093),
    .X(_00928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07193_ (.A0(net3589),
    .A1(net3576),
    .S(net1093),
    .X(_00929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07194_ (.A0(net3576),
    .A1(net3574),
    .S(net1093),
    .X(_00930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07195_ (.A0(net3574),
    .A1(net3556),
    .S(net1093),
    .X(_00931_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07196_ (.A0(net3556),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[4] ),
    .S(net1093),
    .X(_00932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07197_ (.A0(net3654),
    .A1(net1967),
    .S(net1093),
    .X(_00933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07198_ (.A(net1967),
    .B(net1092),
    .Y(_02961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07199_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01409_),
    .A2(net1092),
    .Y(_00934_),
    .B1(_02961_));
 sg13g2_nor2_1 _07200_ (.A(net1935),
    .B(net1091),
    .Y(_02962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07201_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01410_),
    .A2(net1091),
    .Y(_00935_),
    .B1(_02962_));
 sg13g2_nor2_1 _07202_ (.A(net1968),
    .B(net1088),
    .Y(_02963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07203_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01411_),
    .A2(net1088),
    .Y(_00936_),
    .B1(_02963_));
 sg13g2_nand2_1 _07204_ (.Y(_02964_),
    .A(net1933),
    .B(net1088),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07205_ (.B1(_02964_),
    .VDD(VPWR),
    .Y(_00937_),
    .VSS(VGND),
    .A1(_01411_),
    .A2(net1088));
 sg13g2_mux2_1 _07206_ (.A0(net1933),
    .A1(net2105),
    .S(net1089),
    .X(_00938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07207_ (.A(net2105),
    .B(net1088),
    .Y(_02965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07208_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01413_),
    .A2(net1088),
    .Y(_00939_),
    .B1(_02965_));
 sg13g2_nor2_1 _07209_ (.A(net1897),
    .B(net1089),
    .Y(_02966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07210_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01414_),
    .A2(net1089),
    .Y(_00940_),
    .B1(_02966_));
 sg13g2_nor2_1 _07211_ (.A(net1905),
    .B(net1088),
    .Y(_02967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07212_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01415_),
    .A2(net1088),
    .Y(_00941_),
    .B1(_02967_));
 sg13g2_nand2_1 _07213_ (.Y(_02968_),
    .A(net1945),
    .B(net1090),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07214_ (.B1(_02968_),
    .VDD(VPWR),
    .Y(_00942_),
    .VSS(VGND),
    .A1(_01415_),
    .A2(net1089));
 sg13g2_mux2_1 _07215_ (.A0(net1945),
    .A1(net2432),
    .S(net1090),
    .X(_00943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07216_ (.A(net2432),
    .B(net1090),
    .Y(_02969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07217_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01416_),
    .A2(net1090),
    .Y(_00944_),
    .B1(_02969_));
 sg13g2_nor2_1 _07218_ (.A(net1951),
    .B(net1090),
    .Y(_02970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07219_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01417_),
    .A2(net1090),
    .Y(_00945_),
    .B1(_02970_));
 sg13g2_nand2_1 _07220_ (.Y(_02971_),
    .A(net1937),
    .B(net1087),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07221_ (.B1(_02971_),
    .VDD(VPWR),
    .Y(_00946_),
    .VSS(VGND),
    .A1(_01417_),
    .A2(net1086));
 sg13g2_mux2_1 _07222_ (.A0(net1937),
    .A1(net3655),
    .S(net1087),
    .X(_00947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07223_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[19] ),
    .A1(net3644),
    .S(net1086),
    .X(_00948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07224_ (.A0(net3644),
    .A1(net3600),
    .S(net1086),
    .X(_00949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07225_ (.A0(net3600),
    .A1(net3587),
    .S(net1086),
    .X(_00950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07226_ (.A0(net3587),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[23] ),
    .S(net1087),
    .X(_00951_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07227_ (.A0(net3638),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[24] ),
    .S(net1087),
    .X(_00952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07228_ (.A0(net3663),
    .A1(\i_exotiny.i_wb_spi.dat_rx_r[25] ),
    .S(net1086),
    .X(_00953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07229_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[25] ),
    .A1(net3659),
    .S(net1086),
    .X(_00954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07230_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[26] ),
    .A1(net3616),
    .S(net1086),
    .X(_00955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07231_ (.A0(net3616),
    .A1(net3623),
    .S(net1086),
    .X(_00956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07232_ (.A0(net3623),
    .A1(net3646),
    .S(net1092),
    .X(_00957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07233_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[29] ),
    .A1(net3582),
    .S(net1092),
    .X(_00958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07234_ (.A0(\i_exotiny.i_wb_spi.dat_rx_r[30] ),
    .A1(net3530),
    .S(net1092),
    .X(_00959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07235_ (.A(_02518_),
    .B(_02564_),
    .Y(_02972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07236_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1139),
    .A2(_02972_),
    .Y(_02973_),
    .B1(net1166));
 sg13g2_mux2_1 _07237_ (.A0(net3314),
    .A1(net3341),
    .S(net1004),
    .X(_00960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07238_ (.A0(net2889),
    .A1(\i_exotiny._0040_[1] ),
    .S(net1005),
    .X(_00961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07239_ (.A0(net3083),
    .A1(\i_exotiny._0040_[2] ),
    .S(net1004),
    .X(_00962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07240_ (.A0(net2467),
    .A1(net3049),
    .S(net1005),
    .X(_00963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07241_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[8] ),
    .A1(net3314),
    .S(net1007),
    .X(_00964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07242_ (.A0(net2934),
    .A1(net2889),
    .S(net1005),
    .X(_00965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07243_ (.A0(net2361),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[6] ),
    .S(net1003),
    .X(_00966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07244_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[11] ),
    .A1(net2467),
    .S(net1006),
    .X(_00967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07245_ (.A0(net2878),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[8] ),
    .S(net1004),
    .X(_00968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07246_ (.A0(net3089),
    .A1(net2934),
    .S(net1005),
    .X(_00969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07247_ (.A0(net2487),
    .A1(net2361),
    .S(net1003),
    .X(_00970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07248_ (.A0(net3352),
    .A1(net3386),
    .S(net1006),
    .X(_00971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07249_ (.A0(net2311),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[12] ),
    .S(net1004),
    .X(_00972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07250_ (.A0(net2924),
    .A1(net3089),
    .S(net1005),
    .X(_00973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07251_ (.A0(net2339),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[14] ),
    .S(net1003),
    .X(_00974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07252_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[19] ),
    .A1(net3352),
    .S(net1006),
    .X(_00975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07253_ (.A0(net2309),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[16] ),
    .S(net1004),
    .X(_00976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07254_ (.A0(net2713),
    .A1(net2924),
    .S(net1005),
    .X(_00977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07255_ (.A0(net2616),
    .A1(net2339),
    .S(net1003),
    .X(_00978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07256_ (.A0(net2454),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[19] ),
    .S(net1006),
    .X(_00979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07257_ (.A0(net2759),
    .A1(net2309),
    .S(net1004),
    .X(_00980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07258_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[25] ),
    .A1(net2713),
    .S(net1005),
    .X(_00981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07259_ (.A0(net2973),
    .A1(net2616),
    .S(net1003),
    .X(_00982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07260_ (.A0(net2542),
    .A1(net2454),
    .S(net1004),
    .X(_00983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07261_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[28] ),
    .A1(net2759),
    .S(net1003),
    .X(_00984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07262_ (.A0(net2398),
    .A1(net3126),
    .S(net1006),
    .X(_00985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07263_ (.A0(net2614),
    .A1(net2973),
    .S(net1003),
    .X(_00986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07264_ (.A0(net3173),
    .A1(net2542),
    .S(net1006),
    .X(_00987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07265_ (.A0(\i_exotiny._0040_[0] ),
    .A1(net890),
    .S(_02972_),
    .X(_02974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07266_ (.A0(_02974_),
    .A1(net3071),
    .S(net1007),
    .X(_00988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07267_ (.A0(\i_exotiny._0040_[1] ),
    .A1(net883),
    .S(_02972_),
    .X(_02975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07268_ (.A0(_02975_),
    .A1(net2398),
    .S(net1005),
    .X(_00989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07269_ (.A0(\i_exotiny._0040_[2] ),
    .A1(net880),
    .S(_02972_),
    .X(_02976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07270_ (.A0(_02976_),
    .A1(net2614),
    .S(net1003),
    .X(_00990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07271_ (.A0(net3049),
    .A1(net874),
    .S(_02972_),
    .X(_02977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07272_ (.A0(_02977_),
    .A1(net3173),
    .S(net1006),
    .X(_00991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _07273_ (.Y(_02978_),
    .B(_02476_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_02420_));
 sg13g2_o21ai_1 _07274_ (.B1(net1158),
    .VDD(VPWR),
    .Y(_02979_),
    .VSS(VGND),
    .A1(_02423_),
    .A2(_02978_));
 sg13g2_mux2_1 _07275_ (.A0(\i_exotiny._0042_[0] ),
    .A1(net2438),
    .S(net910),
    .X(_00992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07276_ (.A0(net2840),
    .A1(net2654),
    .S(net912),
    .X(_00993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07277_ (.A0(net3168),
    .A1(net3210),
    .S(net912),
    .X(_00994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07278_ (.A0(\i_exotiny._0042_[3] ),
    .A1(net2202),
    .S(net911),
    .X(_00995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07279_ (.A0(net2438),
    .A1(net2767),
    .S(net909),
    .X(_00996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07280_ (.A0(net2654),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[9] ),
    .S(net908),
    .X(_00997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07281_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[6] ),
    .A1(net2584),
    .S(net909),
    .X(_00998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07282_ (.A0(net2202),
    .A1(net2789),
    .S(net911),
    .X(_00999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07283_ (.A0(net2767),
    .A1(net3363),
    .S(net910),
    .X(_01000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07284_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[9] ),
    .A1(net2067),
    .S(net908),
    .X(_01001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07285_ (.A0(net2584),
    .A1(net2907),
    .S(net909),
    .X(_01002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07286_ (.A0(net2789),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[15] ),
    .S(net911),
    .X(_01003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07287_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[12] ),
    .A1(net2715),
    .S(net910),
    .X(_01004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07288_ (.A0(net2067),
    .A1(net2127),
    .S(net908),
    .X(_01005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07289_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[14] ),
    .A1(net2035),
    .S(net909),
    .X(_01006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07290_ (.A0(net2954),
    .A1(net2846),
    .S(net911),
    .X(_01007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07291_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[16] ),
    .A1(net2245),
    .S(net910),
    .X(_01008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07292_ (.A0(net2127),
    .A1(net2295),
    .S(net908),
    .X(_01009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07293_ (.A0(net2035),
    .A1(net3036),
    .S(net909),
    .X(_01010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07294_ (.A0(net2846),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[23] ),
    .S(net911),
    .X(_01011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07295_ (.A0(net2245),
    .A1(net2662),
    .S(net910),
    .X(_01012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07296_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[21] ),
    .A1(net2103),
    .S(net908),
    .X(_01013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07297_ (.A0(net3036),
    .A1(net3059),
    .S(net909),
    .X(_01014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07298_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[23] ),
    .A1(net3471),
    .S(net911),
    .X(_01015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07299_ (.A0(net2662),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[28] ),
    .S(net909),
    .X(_01016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07300_ (.A0(net2103),
    .A1(net2880),
    .S(net908),
    .X(_01017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07301_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[26] ),
    .A1(net2290),
    .S(net908),
    .X(_01018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07302_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[27] ),
    .A1(net2495),
    .S(net911),
    .X(_01019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07303_ (.A0(net890),
    .A1(\i_exotiny._0042_[0] ),
    .S(_02978_),
    .X(_02980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07304_ (.A0(net3232),
    .A1(_02980_),
    .S(net909),
    .X(_01020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07305_ (.A0(net881),
    .A1(net2840),
    .S(_02978_),
    .X(_02981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07306_ (.A0(net2880),
    .A1(_02981_),
    .S(net908),
    .X(_01021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07307_ (.A0(net880),
    .A1(net3168),
    .S(_02978_),
    .X(_02982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07308_ (.A0(net2290),
    .A1(_02982_),
    .S(net912),
    .X(_01022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07309_ (.A0(net872),
    .A1(net3013),
    .S(_02978_),
    .X(_02983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07310_ (.A0(net2495),
    .A1(_02983_),
    .S(net911),
    .X(_01023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07311_ (.Y(_02984_),
    .B(net1212),
    .A_N(net1196),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07312_ (.A0(net1253),
    .A1(net3798),
    .S(net1150),
    .X(_01024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07313_ (.A0(net3690),
    .A1(\i_exotiny._0369_[3] ),
    .S(net1150),
    .X(_01025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07314_ (.A0(net1251),
    .A1(net3768),
    .S(net1151),
    .X(_01026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07315_ (.A0(net1249),
    .A1(net3800),
    .S(net1150),
    .X(_01027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07316_ (.A(net3684),
    .B(net1150),
    .Y(_02985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07317_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01404_),
    .A2(net1151),
    .Y(_01028_),
    .B1(_02985_));
 sg13g2_mux2_1 _07318_ (.A0(net1246),
    .A1(net3759),
    .S(net1150),
    .X(_01029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07319_ (.Y(_02986_),
    .A(net3749),
    .B(net1150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07320_ (.B1(_02986_),
    .VDD(VPWR),
    .Y(_01030_),
    .VSS(VGND),
    .A1(_01382_),
    .A2(net1150));
 sg13g2_nand2_1 _07321_ (.Y(_02987_),
    .A(net3643),
    .B(net1151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07322_ (.B1(_02987_),
    .VDD(VPWR),
    .Y(_01031_),
    .VSS(VGND),
    .A1(_01381_),
    .A2(net1150));
 sg13g2_mux2_1 _07323_ (.A0(net3761),
    .A1(net3457),
    .S(net1151),
    .X(_01032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07324_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1306_ ),
    .A2(_01461_),
    .Y(_02988_),
    .B1(_01598_));
 sg13g2_a21o_2 _07325_ (.A2(_01461_),
    .A1(\i_exotiny._1306_ ),
    .B1(_01598_),
    .X(_02989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07326_ (.A(net1214),
    .B(_02988_),
    .Y(_02990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07327_ (.Y(_02991_),
    .A(net1208),
    .B(_02989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07328_ (.Y(_02992_),
    .A(\i_exotiny._0369_[2] ),
    .B(\i_exotiny._0369_[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07329_ (.Y(_02993_),
    .A(net1214),
    .B(_02992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07330_ (.A(\i_exotiny._0369_[4] ),
    .B(\i_exotiny._0369_[2] ),
    .Y(_02994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07331_ (.Y(_02995_),
    .A(\i_exotiny._0369_[5] ),
    .B(_02994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07332_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[5] ),
    .A2(_02994_),
    .Y(_02996_),
    .B1(\i_exotiny._0369_[20] ));
 sg13g2_nand2_1 _07333_ (.Y(_02997_),
    .A(\i_exotiny._0369_[4] ),
    .B(\i_exotiny._0369_[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07334_ (.Y(_02998_),
    .A(_01404_),
    .B(\i_exotiny._0369_[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07335_ (.Y(_02999_),
    .A(_02997_),
    .B(_02998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07336_ (.Y(_03000_),
    .A(\i_exotiny._0369_[6] ),
    .B(_02994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07337_ (.VDD(VPWR),
    .Y(_03001_),
    .A(_03000_),
    .VSS(VGND));
 sg13g2_nor2_1 _07338_ (.A(_02999_),
    .B(_03001_),
    .Y(_03002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07339_ (.B1(_03002_),
    .VDD(VPWR),
    .Y(_03003_),
    .VSS(VGND),
    .A1(\i_exotiny._0369_[7] ),
    .A2(_02995_));
 sg13g2_nand2_2 _07340_ (.Y(_03004_),
    .A(_02995_),
    .B(_03000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07341_ (.A(_02993_),
    .B(_02996_),
    .C(_03003_),
    .Y(_03005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07342_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3712),
    .A2(net1212),
    .Y(_03006_),
    .B1(_03005_));
 sg13g2_nor2_1 _07343_ (.A(net3739),
    .B(net1078),
    .Y(_03007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07344_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1078),
    .A2(_03006_),
    .Y(_01033_),
    .B1(_03007_));
 sg13g2_and2_1 _07345_ (.A(net2125),
    .B(net1214),
    .X(_03008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07346_ (.B1(_02992_),
    .VDD(VPWR),
    .Y(_03009_),
    .VSS(VGND),
    .A1(_02999_),
    .A2(_03004_));
 sg13g2_a22oi_1 _07347_ (.Y(_03010_),
    .B1(_03008_),
    .B2(_03009_),
    .A2(net1212),
    .A1(net2044),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07348_ (.Y(_03011_),
    .B1(_03004_),
    .B2(_02626_),
    .A2(net1079),
    .A1(net3770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07349_ (.B1(net3771),
    .VDD(VPWR),
    .Y(_01034_),
    .VSS(VGND),
    .A1(net1079),
    .A2(_03010_));
 sg13g2_nor2_1 _07350_ (.A(net3727),
    .B(net1078),
    .Y(_03012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _07351_ (.A(net3307),
    .B_N(_03009_),
    .Y(_03013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07352_ (.A(\i_exotiny._0369_[3] ),
    .B(_02998_),
    .Y(_03014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07353_ (.Y(_03015_),
    .B(_03004_),
    .A_N(net2997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07354_ (.A(net1207),
    .B(_03013_),
    .C(net1148),
    .Y(_03016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07355_ (.Y(_03017_),
    .B1(_03015_),
    .B2(_03016_),
    .A2(net1207),
    .A1(net3010),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07356_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1078),
    .A2(_03017_),
    .Y(_01035_),
    .B1(_03012_));
 sg13g2_and2_1 _07357_ (.A(net2061),
    .B(net1214),
    .X(_03018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07358_ (.Y(_03019_),
    .B1(_03009_),
    .B2(_03018_),
    .A2(net1207),
    .A1(net1949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07359_ (.Y(_03020_),
    .B1(_03004_),
    .B2(_02628_),
    .A2(net1079),
    .A1(net3802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07360_ (.B1(net3803),
    .VDD(VPWR),
    .Y(_01036_),
    .VSS(VGND),
    .A1(net1079),
    .A2(_03019_));
 sg13g2_and2_1 _07361_ (.A(net3647),
    .B(net1213),
    .X(_03021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07362_ (.Y(_03022_),
    .B1(_03009_),
    .B2(_03021_),
    .A2(net1208),
    .A1(net1989),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07363_ (.Y(_03023_),
    .B1(_03004_),
    .B2(_02629_),
    .A2(net1079),
    .A1(net3712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07364_ (.B1(_03023_),
    .VDD(VPWR),
    .Y(_01037_),
    .VSS(VGND),
    .A1(net1079),
    .A2(_03022_));
 sg13g2_nor2_1 _07365_ (.A(net2044),
    .B(_02991_),
    .Y(_03024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07366_ (.Y(_03025_),
    .A(_02992_),
    .B(_02999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07367_ (.A(\i_exotiny._0369_[25] ),
    .B(net1213),
    .X(_03026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07368_ (.Y(_03027_),
    .B1(_03025_),
    .B2(_03026_),
    .A2(net1212),
    .A1(net1996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07369_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1077),
    .A2(_03027_),
    .Y(_01038_),
    .B1(_03024_));
 sg13g2_and2_1 _07370_ (.A(net1872),
    .B(net1217),
    .X(_03028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07371_ (.Y(_03029_),
    .B1(_03025_),
    .B2(_03028_),
    .A2(net1207),
    .A1(net2026),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07372_ (.A(net3010),
    .B(net1078),
    .Y(_03030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07373_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1078),
    .A2(_03029_),
    .Y(_01039_),
    .B1(_03030_));
 sg13g2_nor2_1 _07374_ (.A(net1949),
    .B(net1077),
    .Y(_03031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07375_ (.A(net3584),
    .B(net1213),
    .X(_03032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07376_ (.Y(_03033_),
    .B1(_03025_),
    .B2(_03032_),
    .A2(net1208),
    .A1(\i_exotiny._1160_[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07377_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1077),
    .A2(_03033_),
    .Y(_01040_),
    .B1(_03031_));
 sg13g2_nor2_1 _07378_ (.A(net1989),
    .B(_02991_),
    .Y(_03034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07379_ (.A(\i_exotiny._0369_[28] ),
    .B(net1213),
    .X(_03035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07380_ (.Y(_03036_),
    .B1(_03025_),
    .B2(_03035_),
    .A2(net1210),
    .A1(\i_exotiny._1160_[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07381_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1077),
    .A2(_03036_),
    .Y(_01041_),
    .B1(_03034_));
 sg13g2_and2_1 _07382_ (.A(\i_exotiny._0369_[29] ),
    .B(net1213),
    .X(_03037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07383_ (.Y(_03038_),
    .B1(_03025_),
    .B2(_03037_),
    .A2(net1210),
    .A1(\i_exotiny._1160_[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07384_ (.A(net1996),
    .B(net1077),
    .Y(_03039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07385_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1077),
    .A2(_03038_),
    .Y(_01042_),
    .B1(_03039_));
 sg13g2_nor2_1 _07386_ (.A(net2026),
    .B(net1078),
    .Y(_03040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07387_ (.A(\i_exotiny._0369_[30] ),
    .B(net1214),
    .X(_03041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07388_ (.Y(_03042_),
    .B1(_03025_),
    .B2(_03041_),
    .A2(net1207),
    .A1(\i_exotiny._1160_[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07389_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1078),
    .A2(_03042_),
    .Y(_01043_),
    .B1(_03040_));
 sg13g2_nor2_1 _07390_ (.A(net1955),
    .B(net1077),
    .Y(_03043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07391_ (.A(net3828),
    .B(net1215),
    .X(_03044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07392_ (.Y(_03045_),
    .A(\i_exotiny._0369_[20] ),
    .B(net1214),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07393_ (.Y(_03046_),
    .B1(_03002_),
    .B2(\i_exotiny._1840_[11] ),
    .A2(_03001_),
    .A1(\i_exotiny._0369_[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07394_ (.Y(_03047_),
    .B1(_03046_),
    .B2(_02992_),
    .A2(_03045_),
    .A1(_02993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07395_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._1160_[11] ),
    .A2(net1208),
    .Y(_03048_),
    .B1(_03047_));
 sg13g2_a21oi_1 _07396_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1077),
    .A2(_03048_),
    .Y(_01044_),
    .B1(_03043_));
 sg13g2_nor2_1 _07397_ (.A(\i_exotiny._1160_[12] ),
    .B(net1216),
    .Y(_03049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07398_ (.Y(_03050_),
    .A(_02992_),
    .B(_02998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07399_ (.Y(_03051_),
    .A(\i_exotiny._1840_[11] ),
    .B(_02992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07400_ (.B1(net1214),
    .VDD(VPWR),
    .Y(_03052_),
    .VSS(VGND),
    .A1(_02999_),
    .A2(_03051_));
 sg13g2_a21oi_1 _07401_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[12] ),
    .A2(net1147),
    .Y(_03053_),
    .B1(_03052_));
 sg13g2_nor3_1 _07402_ (.A(net1079),
    .B(_03049_),
    .C(_03053_),
    .Y(_03054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07403_ (.A2(net1079),
    .A1(net2022),
    .B1(_03054_),
    .X(_01045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07404_ (.A(net2010),
    .B(net1216),
    .Y(_03055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07405_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[13] ),
    .A2(net1147),
    .Y(_03056_),
    .B1(_03052_));
 sg13g2_nor3_1 _07406_ (.A(net1085),
    .B(_03055_),
    .C(_03056_),
    .Y(_03057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07407_ (.A2(net1085),
    .A1(net2065),
    .B1(_03057_),
    .X(_01046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07408_ (.A(net2040),
    .B(net1215),
    .Y(_03058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07409_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[14] ),
    .A2(_03050_),
    .Y(_03059_),
    .B1(_03052_));
 sg13g2_nor3_1 _07410_ (.A(net1080),
    .B(_03058_),
    .C(_03059_),
    .Y(_03060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07411_ (.A2(net1080),
    .A1(net2101),
    .B1(_03060_),
    .X(_01047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07412_ (.A(net2020),
    .B(net1215),
    .Y(_03061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07413_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[15] ),
    .A2(net1147),
    .Y(_03062_),
    .B1(_03052_));
 sg13g2_nor3_1 _07414_ (.A(net1083),
    .B(_03061_),
    .C(_03062_),
    .Y(_03063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07415_ (.A2(net1083),
    .A1(net3526),
    .B1(_03063_),
    .X(_01048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07416_ (.A(\i_exotiny._1160_[16] ),
    .B(net1216),
    .Y(_03064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07417_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[16] ),
    .A2(net1147),
    .Y(_03065_),
    .B1(_03052_));
 sg13g2_nor3_1 _07418_ (.A(net1082),
    .B(_03064_),
    .C(_03065_),
    .Y(_03066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07419_ (.A2(net1082),
    .A1(net2077),
    .B1(_03066_),
    .X(_01049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07420_ (.A(\i_exotiny._1160_[17] ),
    .B(net1215),
    .Y(_03067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07421_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[17] ),
    .A2(net1147),
    .Y(_03068_),
    .B1(_03052_));
 sg13g2_nor3_1 _07422_ (.A(net1083),
    .B(_03067_),
    .C(_03068_),
    .Y(_03069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07423_ (.A2(net1082),
    .A1(net2010),
    .B1(_03069_),
    .X(_01050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07424_ (.A(\i_exotiny._1160_[18] ),
    .B(net1215),
    .Y(_03070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07425_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[18] ),
    .A2(net1147),
    .Y(_03071_),
    .B1(_03052_));
 sg13g2_nor3_1 _07426_ (.A(net1081),
    .B(_03070_),
    .C(_03071_),
    .Y(_03072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07427_ (.A2(net1081),
    .A1(net2040),
    .B1(_03072_),
    .X(_01051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07428_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny._0369_[19] ),
    .A2(net1147),
    .Y(_03073_),
    .B1(_03052_));
 sg13g2_nor2_1 _07429_ (.A(\i_exotiny._1160_[19] ),
    .B(net1215),
    .Y(_03074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07430_ (.A(net1081),
    .B(_03073_),
    .C(_03074_),
    .Y(_03075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07431_ (.A2(net1081),
    .A1(net2020),
    .B1(_03075_),
    .X(_01052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07432_ (.A(net3387),
    .B(net1214),
    .X(_03076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07433_ (.A(_03025_),
    .B(_03076_),
    .X(_03077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07434_ (.Y(_03078_),
    .A(_03025_),
    .B(_03076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07435_ (.Y(_03079_),
    .B1(net1148),
    .B2(_03044_),
    .A2(net1209),
    .A1(\i_exotiny._1160_[20] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07436_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3541),
    .A2(net1082),
    .Y(_03080_),
    .B1(_03077_));
 sg13g2_o21ai_1 _07437_ (.B1(_03080_),
    .VDD(VPWR),
    .Y(_01053_),
    .VSS(VGND),
    .A1(net1082),
    .A2(_03079_));
 sg13g2_a22oi_1 _07438_ (.Y(_03081_),
    .B1(_03008_),
    .B2(net1149),
    .A2(net1209),
    .A1(net3535),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07439_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3558),
    .A2(net1082),
    .Y(_03082_),
    .B1(_03077_));
 sg13g2_o21ai_1 _07440_ (.B1(_03082_),
    .VDD(VPWR),
    .Y(_01054_),
    .VSS(VGND),
    .A1(net1083),
    .A2(_03081_));
 sg13g2_and2_1 _07441_ (.A(net3307),
    .B(net1215),
    .X(_03083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07442_ (.Y(_03084_),
    .B1(net1149),
    .B2(_03083_),
    .A2(net1209),
    .A1(\i_exotiny._1160_[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07443_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3565),
    .A2(net1081),
    .Y(_03085_),
    .B1(_03077_));
 sg13g2_o21ai_1 _07444_ (.B1(_03085_),
    .VDD(VPWR),
    .Y(_01055_),
    .VSS(VGND),
    .A1(net1081),
    .A2(_03084_));
 sg13g2_a22oi_1 _07445_ (.Y(_03086_),
    .B1(net1149),
    .B2(_03018_),
    .A2(net1209),
    .A1(net3637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07446_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3686),
    .A2(net1080),
    .Y(_03087_),
    .B1(_03077_));
 sg13g2_o21ai_1 _07447_ (.B1(_03087_),
    .VDD(VPWR),
    .Y(_01056_),
    .VSS(VGND),
    .A1(net1081),
    .A2(_03086_));
 sg13g2_a22oi_1 _07448_ (.Y(_03088_),
    .B1(net1149),
    .B2(_03021_),
    .A2(net1209),
    .A1(net3384),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07449_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3598),
    .A2(net1083),
    .Y(_03089_),
    .B1(_03077_));
 sg13g2_o21ai_1 _07450_ (.B1(_03089_),
    .VDD(VPWR),
    .Y(_01057_),
    .VSS(VGND),
    .A1(net1082),
    .A2(_03088_));
 sg13g2_a22oi_1 _07451_ (.Y(_03090_),
    .B1(net1148),
    .B2(_03026_),
    .A2(net1207),
    .A1(net3360),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07452_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3535),
    .A2(net1080),
    .Y(_03091_),
    .B1(_03077_));
 sg13g2_o21ai_1 _07453_ (.B1(_03091_),
    .VDD(VPWR),
    .Y(_01058_),
    .VSS(VGND),
    .A1(net1082),
    .A2(_03090_));
 sg13g2_a22oi_1 _07454_ (.Y(_03092_),
    .B1(net1148),
    .B2(_03028_),
    .A2(net1207),
    .A1(net3415),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07455_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3609),
    .A2(net1080),
    .Y(_03093_),
    .B1(_03077_));
 sg13g2_o21ai_1 _07456_ (.B1(_03093_),
    .VDD(VPWR),
    .Y(_01059_),
    .VSS(VGND),
    .A1(net1080),
    .A2(_03092_));
 sg13g2_nand2_1 _07457_ (.Y(_03094_),
    .A(net1911),
    .B(net1212),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07458_ (.Y(_03095_),
    .B1(net1148),
    .B2(_03032_),
    .A2(net1208),
    .A1(net1911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07459_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3637),
    .A2(net1080),
    .Y(_03096_),
    .B1(_03077_));
 sg13g2_o21ai_1 _07460_ (.B1(_03096_),
    .VDD(VPWR),
    .Y(_01060_),
    .VSS(VGND),
    .A1(net1080),
    .A2(_03095_));
 sg13g2_nand3_1 _07461_ (.B(net1208),
    .C(_02989_),
    .A(net3384),
    .Y(_03097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07462_ (.Y(_03098_),
    .A(net1148),
    .B(_03035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07463_ (.B(_03097_),
    .C(_03098_),
    .A(_03078_),
    .Y(_01061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07464_ (.B(net1208),
    .C(_02989_),
    .A(net3360),
    .Y(_03099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07465_ (.Y(_03100_),
    .A(net1148),
    .B(_03037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07466_ (.B(_03099_),
    .C(_03100_),
    .A(_03078_),
    .Y(_01062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07467_ (.B(net1207),
    .C(_02989_),
    .A(net3415),
    .Y(_03101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07468_ (.Y(_03102_),
    .A(net1148),
    .B(_03041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07469_ (.B(_03101_),
    .C(_03102_),
    .A(_03078_),
    .Y(_01063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07470_ (.B1(_03076_),
    .VDD(VPWR),
    .Y(_03103_),
    .VSS(VGND),
    .A1(_02997_),
    .A2(net1147));
 sg13g2_o21ai_1 _07471_ (.B1(_03103_),
    .VDD(VPWR),
    .Y(_01064_),
    .VSS(VGND),
    .A1(_02988_),
    .A2(_03094_));
 sg13g2_a21o_1 _07472_ (.A2(net1211),
    .A1(net1241),
    .B1(_03044_),
    .X(_01065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07473_ (.A2(net1211),
    .A1(net1239),
    .B1(_03008_),
    .X(_01066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07474_ (.A2(net1211),
    .A1(net3826),
    .B1(_03083_),
    .X(_01067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07475_ (.A2(net1211),
    .A1(net3825),
    .B1(_03018_),
    .X(_01068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07476_ (.A2(net1211),
    .A1(net3580),
    .B1(_03021_),
    .X(_01069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07477_ (.Y(_03104_),
    .A(_01499_),
    .B(\i_exotiny._1266_ ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07478_ (.Y(_03105_),
    .A(net3819),
    .B(_03104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07479_ (.VDD(VPWR),
    .Y(_03106_),
    .A(net902),
    .VSS(VGND));
 sg13g2_nor2_1 _07480_ (.A(net3820),
    .B(net903),
    .Y(_03107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07481_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01387_),
    .A2(net903),
    .Y(_01070_),
    .B1(_03107_));
 sg13g2_nand2_1 _07482_ (.Y(_03108_),
    .A(net1234),
    .B(net903),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07483_ (.B1(_03108_),
    .VDD(VPWR),
    .Y(_01071_),
    .VSS(VGND),
    .A1(_01393_),
    .A2(net903));
 sg13g2_nand2_1 _07484_ (.Y(_03109_),
    .A(net1233),
    .B(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07485_ (.B1(_03109_),
    .VDD(VPWR),
    .Y(_01072_),
    .VSS(VGND),
    .A1(_01386_),
    .A2(net906));
 sg13g2_nor2_1 _07486_ (.A(net3692),
    .B(net903),
    .Y(_03110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07487_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01390_),
    .A2(net903),
    .Y(_01073_),
    .B1(_03110_));
 sg13g2_nor2_1 _07488_ (.A(net3670),
    .B(net907),
    .Y(_03111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07489_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01391_),
    .A2(net903),
    .Y(_01074_),
    .B1(_03111_));
 sg13g2_nor2_1 _07490_ (.A(net3555),
    .B(net906),
    .Y(_03112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07491_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01393_),
    .A2(net906),
    .Y(_01075_),
    .B1(_03112_));
 sg13g2_nor2_1 _07492_ (.A(net3537),
    .B(net906),
    .Y(_03113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07493_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01386_),
    .A2(net906),
    .Y(_01076_),
    .B1(_03113_));
 sg13g2_mux2_1 _07494_ (.A0(net3626),
    .A1(net3692),
    .S(net907),
    .X(_01077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07495_ (.A0(net3665),
    .A1(net3670),
    .S(net902),
    .X(_01078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07496_ (.A0(net3545),
    .A1(net3555),
    .S(net904),
    .X(_01079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07497_ (.A0(net3547),
    .A1(net3537),
    .S(net905),
    .X(_01080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07498_ (.A0(net3612),
    .A1(net3626),
    .S(net904),
    .X(_01081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07499_ (.A0(net3661),
    .A1(net3665),
    .S(net902),
    .X(_01082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07500_ (.A0(\i_exotiny._0315_[17] ),
    .A1(net3545),
    .S(net904),
    .X(_01083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07501_ (.A0(\i_exotiny._0315_[18] ),
    .A1(net3547),
    .S(net905),
    .X(_01084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07502_ (.A0(\i_exotiny._0315_[19] ),
    .A1(net3612),
    .S(net904),
    .X(_01085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07503_ (.A0(\i_exotiny._0315_[20] ),
    .A1(net3661),
    .S(net901),
    .X(_01086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07504_ (.A0(net3318),
    .A1(net3706),
    .S(net902),
    .X(_01087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07505_ (.A0(\i_exotiny._0315_[22] ),
    .A1(net3549),
    .S(net905),
    .X(_01088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07506_ (.A0(net3185),
    .A1(net3625),
    .S(net904),
    .X(_01089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07507_ (.A0(net2841),
    .A1(\i_exotiny._0315_[20] ),
    .S(net901),
    .X(_01090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07508_ (.A0(net3220),
    .A1(net3318),
    .S(net902),
    .X(_01091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07509_ (.A0(net3113),
    .A1(\i_exotiny._0315_[22] ),
    .S(net905),
    .X(_01092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07510_ (.A0(net3052),
    .A1(net3185),
    .S(net904),
    .X(_01093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07511_ (.A0(net2099),
    .A1(net2841),
    .S(net901),
    .X(_01094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07512_ (.A0(\i_exotiny._0315_[29] ),
    .A1(net3220),
    .S(net901),
    .X(_01095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07513_ (.A0(net3377),
    .A1(net3113),
    .S(net904),
    .X(_01096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07514_ (.A0(net2024),
    .A1(net3052),
    .S(net904),
    .X(_01097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07515_ (.Y(_03114_),
    .A(net2099),
    .B(net901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07516_ (.A(_01499_),
    .B(_02437_),
    .Y(_03115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07517_ (.B1(_03106_),
    .VDD(VPWR),
    .Y(_03116_),
    .VSS(VGND),
    .A1(_01500_),
    .A2(_02014_));
 sg13g2_o21ai_1 _07518_ (.B1(_03114_),
    .VDD(VPWR),
    .Y(_01098_),
    .VSS(VGND),
    .A1(_03115_),
    .A2(_03116_));
 sg13g2_a21o_1 _07519_ (.A2(_01945_),
    .A1(_01499_),
    .B1(net901),
    .X(_03117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07520_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01500_),
    .A2(_02453_),
    .Y(_03118_),
    .B1(_03117_));
 sg13g2_a21o_1 _07521_ (.A2(net901),
    .A1(net3570),
    .B1(_03118_),
    .X(_01099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07522_ (.Y(_03119_),
    .A(net3377),
    .B(net902),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07523_ (.A(net3470),
    .B(_02462_),
    .Y(_03120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07524_ (.B1(_03106_),
    .VDD(VPWR),
    .Y(_03121_),
    .VSS(VGND),
    .A1(_01500_),
    .A2(_01872_));
 sg13g2_o21ai_1 _07525_ (.B1(_03119_),
    .VDD(VPWR),
    .Y(_01100_),
    .VSS(VGND),
    .A1(_03120_),
    .A2(_03121_));
 sg13g2_nand2_1 _07526_ (.Y(_03122_),
    .A(net2024),
    .B(net901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07527_ (.A(_01499_),
    .B(_02471_),
    .Y(_03123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _07528_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01814_),
    .C1(_01500_),
    .B1(_01752_),
    .A1(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ),
    .Y(_03124_),
    .A2(_01686_));
 sg13g2_nand2b_1 _07529_ (.Y(_03125_),
    .B(_03106_),
    .A_N(_03124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07530_ (.B1(_03122_),
    .VDD(VPWR),
    .Y(_01101_),
    .VSS(VGND),
    .A1(_03123_),
    .A2(_03125_));
 sg13g2_nor4_2 _07531_ (.A(net1270),
    .B(net1273),
    .C(net3694),
    .Y(_03126_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1893));
 sg13g2_nand2_1 _07532_ (.Y(_03127_),
    .A(_01363_),
    .B(_03126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07533_ (.B(\i_exotiny._1265_ ),
    .C(_01474_),
    .A(net3819),
    .Y(_03128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07534_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03127_),
    .A2(_03128_),
    .Y(_01102_),
    .B1(net1196));
 sg13g2_or2_1 _07535_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_03129_),
    .B(net3824),
    .A(net3832));
 sg13g2_nand3_1 _07536_ (.B(_03126_),
    .C(_03129_),
    .A(_01442_),
    .Y(_03130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07537_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03128_),
    .A2(_03130_),
    .Y(_01103_),
    .B1(net1196));
 sg13g2_nand2_1 _07538_ (.Y(_03131_),
    .A(_01362_),
    .B(_01442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07539_ (.B(_03126_),
    .C(_03131_),
    .A(_01443_),
    .Y(_03132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07540_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03128_),
    .A2(_03132_),
    .Y(_01104_),
    .B1(net1196));
 sg13g2_nand2_2 _07541_ (.Y(_03133_),
    .A(net3466),
    .B(net1290),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07542_ (.VDD(VPWR),
    .Y(_03134_),
    .A(_03133_),
    .VSS(VGND));
 sg13g2_nor2_1 _07543_ (.A(net1883),
    .B(_03133_),
    .Y(_01105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07544_ (.Y(_03135_),
    .A(net1883),
    .B(net3586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07545_ (.A(_03133_),
    .B(_03135_),
    .Y(_01106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07546_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1883),
    .A2(\i_exotiny.i_rstctl.cnt[1] ),
    .Y(_03136_),
    .B1(net2298));
 sg13g2_and3_1 _07547_ (.X(_03137_),
    .A(net1883),
    .B(net3586),
    .C(net2298),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07548_ (.A(_03133_),
    .B(net2299),
    .C(_03137_),
    .Y(_01107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07549_ (.A(net3658),
    .B(_03137_),
    .Y(_03138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07550_ (.A(net3658),
    .B(_03137_),
    .X(_03139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07551_ (.A(_03133_),
    .B(_03138_),
    .C(_03139_),
    .Y(_01108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07552_ (.A(net3763),
    .B(_03139_),
    .X(_03140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07553_ (.B1(_03134_),
    .VDD(VPWR),
    .Y(_03141_),
    .VSS(VGND),
    .A1(net3763),
    .A2(_03139_));
 sg13g2_nor2_1 _07554_ (.A(_03140_),
    .B(_03141_),
    .Y(_01109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07555_ (.A(net3681),
    .B(_03140_),
    .X(_03142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07556_ (.B1(_03134_),
    .VDD(VPWR),
    .Y(_03143_),
    .VSS(VGND),
    .A1(net3681),
    .A2(_03140_));
 sg13g2_nor2_1 _07557_ (.A(_03142_),
    .B(_03143_),
    .Y(_01110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07558_ (.B1(_03134_),
    .VDD(VPWR),
    .Y(_03144_),
    .VSS(VGND),
    .A1(net1970),
    .A2(_03142_));
 sg13g2_a21oi_1 _07559_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1970),
    .A2(_03142_),
    .Y(_01111_),
    .B1(_03144_));
 sg13g2_nor4_1 _07560_ (.A(net3833),
    .B(net3520),
    .C(net3724),
    .D(_01521_),
    .Y(_03145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07561_ (.A(net1225),
    .B(net1231),
    .C(_03145_),
    .Y(_01112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07562_ (.A(net3520),
    .B(net3724),
    .C(_02178_),
    .Y(_03146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _07563_ (.A(net3520),
    .B(_01527_),
    .C(_02177_),
    .D(_03146_),
    .Y(_03147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07564_ (.A(net3699),
    .B(net1231),
    .Y(_03148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07565_ (.Y(_03149_),
    .A(net1283),
    .B(_01486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07566_ (.A(_03147_),
    .B(_03148_),
    .C(_03149_),
    .Y(_01113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07567_ (.A2(_01493_),
    .A1(net3520),
    .B1(_03146_),
    .X(_03150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _07568_ (.A(\i_exotiny._1737_ ),
    .B(_01527_),
    .C(_01545_),
    .D(_03150_),
    .Y(_03151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07569_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3699),
    .A2(net1231),
    .Y(_03152_),
    .B1(\i_exotiny.i_wb_qspi_mem.cnt_r[2] ));
 sg13g2_nor4_1 _07570_ (.A(net1225),
    .B(_01487_),
    .C(_03151_),
    .D(net3700),
    .Y(_01114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07571_ (.A(net1830),
    .B(net1204),
    .Y(_01115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07572_ (.A(net3201),
    .B(net1830),
    .Y(_03153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07573_ (.A(net3201),
    .B(net1830),
    .X(_03154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07574_ (.A(net1204),
    .B(_03153_),
    .C(_03154_),
    .Y(_01116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07575_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net3756),
    .A2(_03154_),
    .Y(_03155_),
    .B1(net1204));
 sg13g2_o21ai_1 _07576_ (.B1(_03155_),
    .VDD(VPWR),
    .Y(_03156_),
    .VSS(VGND),
    .A1(net3756),
    .A2(_03154_));
 sg13g2_inv_1 _07577_ (.VDD(VPWR),
    .Y(_01117_),
    .A(_03156_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07578_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_wdg_top.clk_div_inst.cnt[2] ),
    .A2(_03154_),
    .Y(_03157_),
    .B1(net1885));
 sg13g2_and3_1 _07579_ (.X(_03158_),
    .A(net3844),
    .B(net1885),
    .C(_03154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07580_ (.A(net1204),
    .B(net1886),
    .C(_03158_),
    .Y(_01118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07581_ (.A(net3627),
    .B(_03158_),
    .X(_03159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07582_ (.B1(net1179),
    .VDD(VPWR),
    .Y(_03160_),
    .VSS(VGND),
    .A1(net3627),
    .A2(_03158_));
 sg13g2_nor2_1 _07583_ (.A(_03159_),
    .B(net3628),
    .Y(_01119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07584_ (.Y(_03161_),
    .A(net3671),
    .B(_03159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07585_ (.A(net1204),
    .B(_03161_),
    .Y(_01120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07586_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_wdg_top.clk_div_inst.cnt[5] ),
    .A2(_03159_),
    .Y(_03162_),
    .B1(net1913));
 sg13g2_and3_1 _07587_ (.X(_03163_),
    .A(net3843),
    .B(net1913),
    .C(_03159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07588_ (.A(net1204),
    .B(net1914),
    .C(_03163_),
    .Y(_01121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07589_ (.A(net2028),
    .B(_03163_),
    .Y(_03164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07590_ (.A(net2028),
    .B(_03163_),
    .X(_03165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07591_ (.A(net1206),
    .B(net2029),
    .C(_03165_),
    .Y(_01122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07592_ (.A(net3642),
    .B(_03165_),
    .X(_03166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07593_ (.B1(net1179),
    .VDD(VPWR),
    .Y(_03167_),
    .VSS(VGND),
    .A1(net3642),
    .A2(_03165_));
 sg13g2_nor2_1 _07594_ (.A(_03166_),
    .B(_03167_),
    .Y(_01123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07595_ (.Y(_03168_),
    .A(net3607),
    .B(_03166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07596_ (.A(net1205),
    .B(net3608),
    .Y(_01124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07597_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_wdg_top.clk_div_inst.cnt[9] ),
    .A2(_03166_),
    .Y(_03169_),
    .B1(net1877));
 sg13g2_and3_2 _07598_ (.X(_03170_),
    .A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[9] ),
    .B(net1877),
    .C(_03166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07599_ (.A(net1205),
    .B(net1878),
    .C(_03170_),
    .Y(_01125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07600_ (.Y(_03171_),
    .A(net3578),
    .B(_03170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07601_ (.A(net1205),
    .B(net3579),
    .Y(_01126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07602_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_wdg_top.clk_div_inst.cnt[11] ),
    .A2(_03170_),
    .Y(_03172_),
    .B1(net1890));
 sg13g2_and3_1 _07603_ (.X(_03173_),
    .A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[11] ),
    .B(net1890),
    .C(_03170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07604_ (.A(net1206),
    .B(net1891),
    .C(_03173_),
    .Y(_01127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07605_ (.A(net3235),
    .B(_03173_),
    .Y(_03174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07606_ (.A(net3235),
    .B(_03173_),
    .X(_03175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07607_ (.A(net1205),
    .B(net3236),
    .C(_03175_),
    .Y(_01128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07608_ (.A(net3722),
    .B(_03175_),
    .X(_03176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07609_ (.B1(\i_exotiny._0000_ ),
    .VDD(VPWR),
    .Y(_03177_),
    .VSS(VGND),
    .A1(net3722),
    .A2(_03175_));
 sg13g2_nor2_1 _07610_ (.A(_03176_),
    .B(net3723),
    .Y(_01129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07611_ (.Y(_03178_),
    .A(net3649),
    .B(_03176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07612_ (.A(net1205),
    .B(net3650),
    .Y(_01130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07613_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\i_exotiny.i_wdg_top.clk_div_inst.cnt[15] ),
    .A2(_03176_),
    .Y(_03179_),
    .B1(net1880));
 sg13g2_and3_1 _07614_ (.X(_03180_),
    .A(net3842),
    .B(net1880),
    .C(_03176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07615_ (.A(net1205),
    .B(net1881),
    .C(_03180_),
    .Y(_01131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07616_ (.A(net2054),
    .B(_03180_),
    .Y(_03181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07617_ (.A(net2054),
    .B(_03180_),
    .X(_03182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07618_ (.A(net1205),
    .B(net2055),
    .C(_03182_),
    .Y(_01132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07619_ (.A(net3569),
    .B(_03182_),
    .X(_03183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07620_ (.B1(\i_exotiny._0000_ ),
    .VDD(VPWR),
    .Y(_03184_),
    .VSS(VGND),
    .A1(net3569),
    .A2(_03182_));
 sg13g2_nor2_1 _07621_ (.A(_03183_),
    .B(_03184_),
    .Y(_01133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07622_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1228),
    .A2(_03183_),
    .Y(_03185_),
    .B1(net1205));
 sg13g2_o21ai_1 _07623_ (.B1(_03185_),
    .VDD(VPWR),
    .Y(_03186_),
    .VSS(VGND),
    .A1(net1228),
    .A2(_03183_));
 sg13g2_inv_1 _07624_ (.VDD(VPWR),
    .Y(_01134_),
    .A(_03186_),
    .VSS(VGND));
 sg13g2_nor2_2 _07625_ (.A(_02477_),
    .B(_02517_),
    .Y(_03187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _07626_ (.A2(_03187_),
    .A1(net1141),
    .B1(net1168),
    .X(_03188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07627_ (.A0(\i_exotiny._0024_[0] ),
    .A1(net3105),
    .S(net899),
    .X(_01135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07628_ (.A0(\i_exotiny._0024_[1] ),
    .A1(net2186),
    .S(net898),
    .X(_01136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07629_ (.A0(\i_exotiny._0024_[2] ),
    .A1(net2462),
    .S(net897),
    .X(_01137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07630_ (.A0(\i_exotiny._0024_[3] ),
    .A1(net2917),
    .S(net896),
    .X(_01138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07631_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[4] ),
    .A1(net2097),
    .S(net899),
    .X(_01139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07632_ (.A0(net2186),
    .A1(net2607),
    .S(net898),
    .X(_01140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07633_ (.A0(net2462),
    .A1(net2686),
    .S(net897),
    .X(_01141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07634_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[7] ),
    .A1(net2859),
    .S(net896),
    .X(_01142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07635_ (.A0(net2097),
    .A1(net2958),
    .S(net899),
    .X(_01143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07636_ (.A0(net2607),
    .A1(net3190),
    .S(net898),
    .X(_01144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07637_ (.A0(net2686),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[14] ),
    .S(net897),
    .X(_01145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07638_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[11] ),
    .A1(net2706),
    .S(net896),
    .X(_01146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07639_ (.A0(net2958),
    .A1(net2785),
    .S(net899),
    .X(_01147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07640_ (.A0(net3190),
    .A1(net3311),
    .S(net898),
    .X(_01148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07641_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[14] ),
    .A1(net3338),
    .S(net897),
    .X(_01149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07642_ (.A0(net2706),
    .A1(net2952),
    .S(net896),
    .X(_01150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07643_ (.A0(net2785),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[20] ),
    .S(net899),
    .X(_01151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07644_ (.A0(net3311),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[21] ),
    .S(net898),
    .X(_01152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07645_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[18] ),
    .A1(net2130),
    .S(net897),
    .X(_01153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07646_ (.A0(net2952),
    .A1(net3070),
    .S(net896),
    .X(_01154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07647_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[20] ),
    .A1(net2236),
    .S(net899),
    .X(_01155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07648_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[21] ),
    .A1(net2396),
    .S(net898),
    .X(_01156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07649_ (.A0(net2130),
    .A1(net3004),
    .S(net900),
    .X(_01157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07650_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[23] ),
    .A1(net2349),
    .S(net896),
    .X(_01158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07651_ (.A0(net2236),
    .A1(net3085),
    .S(net899),
    .X(_01159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07652_ (.A0(net2396),
    .A1(net2888),
    .S(net898),
    .X(_01160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07653_ (.A0(net3004),
    .A1(net2296),
    .S(net897),
    .X(_01161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07654_ (.A0(net2349),
    .A1(net3145),
    .S(net896),
    .X(_01162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07655_ (.A0(\i_exotiny._0024_[0] ),
    .A1(net889),
    .S(_03187_),
    .X(_03189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07656_ (.A0(net3085),
    .A1(_03189_),
    .S(net899),
    .X(_01163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07657_ (.A0(net3006),
    .A1(net882),
    .S(_03187_),
    .X(_03190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07658_ (.A0(net2888),
    .A1(_03190_),
    .S(net898),
    .X(_01164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07659_ (.A0(\i_exotiny._0024_[2] ),
    .A1(net879),
    .S(_03187_),
    .X(_03191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07660_ (.A0(net2296),
    .A1(_03191_),
    .S(net896),
    .X(_01165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07661_ (.A0(\i_exotiny._0024_[3] ),
    .A1(net873),
    .S(_03187_),
    .X(_03192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07662_ (.A0(net3145),
    .A1(_03192_),
    .S(net897),
    .X(_01166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07663_ (.A(_02492_),
    .B(_02532_),
    .Y(_03193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _07664_ (.A2(_03193_),
    .A1(net1138),
    .B1(net1165),
    .X(_03194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07665_ (.A0(\i_exotiny._0030_[0] ),
    .A1(net2182),
    .S(net1000),
    .X(_01167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07666_ (.A0(net3319),
    .A1(net2535),
    .S(net999),
    .X(_01168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07667_ (.A0(net2511),
    .A1(net2899),
    .S(net1001),
    .X(_01169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07668_ (.A0(\i_exotiny._0030_[3] ),
    .A1(net2633),
    .S(net1001),
    .X(_01170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07669_ (.A0(net2182),
    .A1(net2980),
    .S(net1000),
    .X(_01171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07670_ (.A0(net2535),
    .A1(net2301),
    .S(net998),
    .X(_01172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07671_ (.A0(net2899),
    .A1(net3062),
    .S(net1001),
    .X(_01173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07672_ (.A0(net2633),
    .A1(net2882),
    .S(net1001),
    .X(_01174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07673_ (.A0(net2980),
    .A1(net3163),
    .S(net1002),
    .X(_01175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07674_ (.A0(net2301),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[13] ),
    .S(net998),
    .X(_01176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07675_ (.A0(net3062),
    .A1(net3434),
    .S(net1002),
    .X(_01177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07676_ (.A0(net2882),
    .A1(net2960),
    .S(net1001),
    .X(_01178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07677_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[12] ),
    .A1(net2420),
    .S(net1002),
    .X(_01179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07678_ (.A0(net3138),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[17] ),
    .S(net998),
    .X(_01180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07679_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[14] ),
    .A1(net3181),
    .S(net1001),
    .X(_01181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07680_ (.A0(net2960),
    .A1(net3196),
    .S(net998),
    .X(_01182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07681_ (.A0(net2420),
    .A1(net3238),
    .S(net1000),
    .X(_01183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07682_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[17] ),
    .A1(net2194),
    .S(net998),
    .X(_01184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07683_ (.A0(net3181),
    .A1(net2499),
    .S(net1001),
    .X(_01185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07684_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[19] ),
    .A1(net2176),
    .S(net998),
    .X(_01186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07685_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[20] ),
    .A1(net2526),
    .S(net1000),
    .X(_01187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07686_ (.A0(net2194),
    .A1(net2978),
    .S(net998),
    .X(_01188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07687_ (.A0(net2499),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[26] ),
    .S(net1001),
    .X(_01189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07688_ (.A0(net2176),
    .A1(net2974),
    .S(net999),
    .X(_01190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07689_ (.A0(net2526),
    .A1(net2976),
    .S(net1000),
    .X(_01191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07690_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[25] ),
    .A1(net2727),
    .S(net999),
    .X(_01192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07691_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[26] ),
    .A1(net2172),
    .S(net1000),
    .X(_01193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07692_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[27] ),
    .A1(net2209),
    .S(net999),
    .X(_01194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07693_ (.A0(\i_exotiny._0030_[0] ),
    .A1(net887),
    .S(_03193_),
    .X(_03195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07694_ (.A0(net2976),
    .A1(_03195_),
    .S(net1000),
    .X(_01195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07695_ (.A0(net3319),
    .A1(net882),
    .S(_03193_),
    .X(_03196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07696_ (.A0(net2727),
    .A1(_03196_),
    .S(net999),
    .X(_01196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07697_ (.A0(net2511),
    .A1(net877),
    .S(_03193_),
    .X(_03197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07698_ (.A0(net2172),
    .A1(_03197_),
    .S(net1000),
    .X(_01197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07699_ (.A0(net3009),
    .A1(net873),
    .S(_03193_),
    .X(_03198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07700_ (.A0(net2209),
    .A1(_03198_),
    .S(net998),
    .X(_01198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07701_ (.A(_02419_),
    .B(_02477_),
    .Y(_03199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07702_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1142),
    .A2(_03199_),
    .Y(_03200_),
    .B1(net1163));
 sg13g2_mux2_1 _07703_ (.A0(net2992),
    .A1(\i_exotiny._0027_[0] ),
    .S(net994),
    .X(_01199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07704_ (.A0(net2959),
    .A1(net3075),
    .S(net996),
    .X(_01200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07705_ (.A0(net2724),
    .A1(net2613),
    .S(net996),
    .X(_01201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07706_ (.A0(net3490),
    .A1(net3459),
    .S(net996),
    .X(_01202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07707_ (.A0(net2990),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[4] ),
    .S(net994),
    .X(_01203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07708_ (.A0(net2545),
    .A1(net2959),
    .S(net994),
    .X(_01204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07709_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[10] ),
    .A1(net2724),
    .S(net996),
    .X(_01205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07710_ (.A0(net3176),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[7] ),
    .S(net995),
    .X(_01206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07711_ (.A0(net2335),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[8] ),
    .S(net993),
    .X(_01207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07712_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[13] ),
    .A1(net2545),
    .S(net997),
    .X(_01208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07713_ (.A0(net3271),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[10] ),
    .S(net995),
    .X(_01209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07714_ (.A0(net3198),
    .A1(net3176),
    .S(net995),
    .X(_01210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07715_ (.A0(net2916),
    .A1(net2335),
    .S(net993),
    .X(_01211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07716_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[17] ),
    .A1(net2579),
    .S(net994),
    .X(_01212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07717_ (.A0(net2422),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[14] ),
    .S(net995),
    .X(_01213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07718_ (.A0(net2568),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[15] ),
    .S(net995),
    .X(_01214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07719_ (.A0(net3090),
    .A1(net2916),
    .S(net993),
    .X(_01215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07720_ (.A0(net2748),
    .A1(net3079),
    .S(net994),
    .X(_01216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07721_ (.A0(net2642),
    .A1(net2422),
    .S(net995),
    .X(_01217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07722_ (.A0(net2885),
    .A1(net2568),
    .S(net995),
    .X(_01218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07723_ (.A0(net2048),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[20] ),
    .S(net993),
    .X(_01219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07724_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[25] ),
    .A1(net2748),
    .S(net993),
    .X(_01220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07725_ (.A0(net3453),
    .A1(net2642),
    .S(net996),
    .X(_01221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07726_ (.A0(net2387),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[23] ),
    .S(net993),
    .X(_01222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07727_ (.A0(net2839),
    .A1(net2048),
    .S(net993),
    .X(_01223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07728_ (.A0(net2379),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[25] ),
    .S(net997),
    .X(_01224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07729_ (.A0(net2517),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[26] ),
    .S(net995),
    .X(_01225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07730_ (.A0(net2547),
    .A1(net2387),
    .S(net993),
    .X(_01226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07731_ (.A0(net3294),
    .A1(net886),
    .S(_03199_),
    .X(_03201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07732_ (.A0(_03201_),
    .A1(net2839),
    .S(net994),
    .X(_01227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07733_ (.A0(net3075),
    .A1(net881),
    .S(_03199_),
    .X(_03202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07734_ (.A0(_03202_),
    .A1(net2379),
    .S(net994),
    .X(_01228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07735_ (.A0(net2613),
    .A1(net876),
    .S(_03199_),
    .X(_03203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07736_ (.A0(_03203_),
    .A1(net2517),
    .S(net996),
    .X(_01229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07737_ (.A0(net3459),
    .A1(net872),
    .S(_03199_),
    .X(_03204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07738_ (.A0(_03204_),
    .A1(net2547),
    .S(net996),
    .X(_01230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07739_ (.A(net1227),
    .B(_01576_),
    .C(net1118),
    .Y(_03205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07740_ (.A(net1119),
    .B(_02946_),
    .Y(_03206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07741_ (.Y(_03207_),
    .A(net3805),
    .B(_03206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07742_ (.B1(_03207_),
    .VDD(VPWR),
    .Y(_03208_),
    .VSS(VGND),
    .A1(net2106),
    .A2(_03206_));
 sg13g2_xnor2_1 _07743_ (.Y(_01231_),
    .A(_03205_),
    .B(_03208_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07744_ (.B(net1116),
    .C(net1060),
    .A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data [0]),
    .Y(_03209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07745_ (.B1(_03209_),
    .VDD(VPWR),
    .Y(_01232_),
    .VSS(VGND),
    .A1(_01397_),
    .A2(net1060));
 sg13g2_nor2_2 _07746_ (.A(_02477_),
    .B(_02564_),
    .Y(_03210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _07747_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(net1166),
    .Y(_03211_),
    .A2(_03210_),
    .A1(net1139));
 sg13g2_mux2_1 _07748_ (.A0(net3157),
    .A1(\i_exotiny._0026_[0] ),
    .S(net991),
    .X(_01233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07749_ (.A0(net2600),
    .A1(\i_exotiny._0026_[1] ),
    .S(net989),
    .X(_01234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07750_ (.A0(net3256),
    .A1(net3270),
    .S(net989),
    .X(_01235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07751_ (.A0(net2460),
    .A1(net2964),
    .S(net988),
    .X(_01236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07752_ (.A0(net3224),
    .A1(net3157),
    .S(net991),
    .X(_01237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07753_ (.A0(net2900),
    .A1(net2600),
    .S(net991),
    .X(_01238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07754_ (.A0(net3057),
    .A1(net3256),
    .S(net988),
    .X(_01239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07755_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[11] ),
    .A1(net2460),
    .S(net990),
    .X(_01240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07756_ (.A0(net2404),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[8] ),
    .S(net991),
    .X(_01241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07757_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[13] ),
    .A1(net2900),
    .S(net991),
    .X(_01242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07758_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[14] ),
    .A1(net3057),
    .S(net988),
    .X(_01243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07759_ (.A0(net2743),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[11] ),
    .S(net990),
    .X(_01244_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07760_ (.A0(net3170),
    .A1(net2404),
    .S(net991),
    .X(_01245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07761_ (.A0(net2241),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[13] ),
    .S(net992),
    .X(_01246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07762_ (.A0(net2581),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[14] ),
    .S(net988),
    .X(_01247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07763_ (.A0(net2780),
    .A1(net2743),
    .S(net990),
    .X(_01248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07764_ (.A0(net2837),
    .A1(net3170),
    .S(net992),
    .X(_01249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07765_ (.A0(net2951),
    .A1(net2241),
    .S(net992),
    .X(_01250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07766_ (.A0(net3317),
    .A1(net2581),
    .S(net989),
    .X(_01251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07767_ (.A0(net2519),
    .A1(net2780),
    .S(net990),
    .X(_01252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07768_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[24] ),
    .A1(net2837),
    .S(net992),
    .X(_01253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07769_ (.A0(net2696),
    .A1(net2951),
    .S(net991),
    .X(_01254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07770_ (.A0(net2132),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[22] ),
    .S(net988),
    .X(_01255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07771_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[27] ),
    .A1(net2519),
    .S(net990),
    .X(_01256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07772_ (.A0(net3007),
    .A1(net3290),
    .S(net990),
    .X(_01257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07773_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[29] ),
    .A1(net2696),
    .S(net991),
    .X(_01258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07774_ (.A0(net3321),
    .A1(net2132),
    .S(net988),
    .X(_01259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07775_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[31] ),
    .A1(net2559),
    .S(net990),
    .X(_01260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07776_ (.A0(\i_exotiny._0026_[0] ),
    .A1(net888),
    .S(_03210_),
    .X(_03212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07777_ (.A0(_03212_),
    .A1(net3007),
    .S(net990),
    .X(_01261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07778_ (.A0(\i_exotiny._0026_[1] ),
    .A1(net883),
    .S(_03210_),
    .X(_03213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07779_ (.A0(_03213_),
    .A1(net3050),
    .S(net989),
    .X(_01262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07780_ (.A0(net3270),
    .A1(net878),
    .S(_03210_),
    .X(_03214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07781_ (.A0(_03214_),
    .A1(net3321),
    .S(net988),
    .X(_01263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07782_ (.A0(\i_exotiny._0026_[3] ),
    .A1(net874),
    .S(_03210_),
    .X(_03215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07783_ (.A0(_03215_),
    .A1(net2853),
    .S(net988),
    .X(_01264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07784_ (.A(_02485_),
    .B(_02518_),
    .Y(_03216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _07785_ (.A2(_03216_),
    .A1(net1138),
    .B1(net1165),
    .X(_03217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07786_ (.A0(\i_exotiny._0023_[0] ),
    .A1(net3227),
    .S(net894),
    .X(_01265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07787_ (.A0(\i_exotiny._0023_[1] ),
    .A1(net3203),
    .S(net895),
    .X(_01266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07788_ (.A0(net3525),
    .A1(net3481),
    .S(net892),
    .X(_01267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07789_ (.A0(net3249),
    .A1(net3508),
    .S(net892),
    .X(_01268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07790_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[4] ),
    .A1(net2071),
    .S(net893),
    .X(_01269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07791_ (.A0(net3203),
    .A1(net2833),
    .S(net894),
    .X(_01270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07792_ (.A0(net3481),
    .A1(net3323),
    .S(net894),
    .X(_01271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07793_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[7] ),
    .A1(net3292),
    .S(net891),
    .X(_01272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07794_ (.A0(net2071),
    .A1(net2935),
    .S(net893),
    .X(_01273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07795_ (.A0(net2833),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[13] ),
    .S(net894),
    .X(_01274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07796_ (.A0(net3323),
    .A1(net2751),
    .S(net893),
    .X(_01275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07797_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[11] ),
    .A1(net2251),
    .S(net891),
    .X(_01276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07798_ (.A0(net2935),
    .A1(net2869),
    .S(net893),
    .X(_01277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07799_ (.A0(net3340),
    .A1(net2625),
    .S(net894),
    .X(_01278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07800_ (.A0(net2751),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[18] ),
    .S(net893),
    .X(_01279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07801_ (.A0(net2251),
    .A1(net3108),
    .S(net891),
    .X(_01280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07802_ (.A0(net2869),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[20] ),
    .S(net893),
    .X(_01281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07803_ (.A0(net2625),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[21] ),
    .S(net894),
    .X(_01282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07804_ (.A0(net3218),
    .A1(net2862),
    .S(net892),
    .X(_01283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07805_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[19] ),
    .A1(net2345),
    .S(net891),
    .X(_01284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07806_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[20] ),
    .A1(net3225),
    .S(net895),
    .X(_01285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07807_ (.A0(net2850),
    .A1(net2680),
    .S(net894),
    .X(_01286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07808_ (.A0(net2862),
    .A1(net2733),
    .S(net892),
    .X(_01287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07809_ (.A0(net2345),
    .A1(net2781),
    .S(net891),
    .X(_01288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07810_ (.A0(net3225),
    .A1(net3017),
    .S(net893),
    .X(_01289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07811_ (.A0(net2680),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[29] ),
    .S(net894),
    .X(_01290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07812_ (.A0(net2733),
    .A1(net2704),
    .S(net891),
    .X(_01291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07813_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[27] ),
    .A1(net2497),
    .S(net891),
    .X(_01292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07814_ (.A0(\i_exotiny._0023_[0] ),
    .A1(net887),
    .S(_03216_),
    .X(_03218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07815_ (.A0(net3017),
    .A1(_03218_),
    .S(net893),
    .X(_01293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07816_ (.A0(\i_exotiny._0023_[1] ),
    .A1(net884),
    .S(_03216_),
    .X(_03219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07817_ (.A0(net3375),
    .A1(_03219_),
    .S(net892),
    .X(_01294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07818_ (.A0(\i_exotiny._0023_[2] ),
    .A1(net879),
    .S(_03216_),
    .X(_03220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07819_ (.A0(net2704),
    .A1(_03220_),
    .S(net892),
    .X(_01295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07820_ (.A0(net3249),
    .A1(net875),
    .S(_03216_),
    .X(_03221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07821_ (.A0(net2497),
    .A1(_03221_),
    .S(net891),
    .X(_01296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07822_ (.A(_02477_),
    .B(_02525_),
    .Y(_03222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1138),
    .A2(_03222_),
    .Y(_03223_),
    .B1(net1168));
 sg13g2_mux2_1 _07824_ (.A0(net2134),
    .A1(\i_exotiny._0022_[0] ),
    .S(net987),
    .X(_01297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07825_ (.A0(net3491),
    .A1(\i_exotiny._0022_[1] ),
    .S(net985),
    .X(_01298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07826_ (.A0(net2162),
    .A1(\i_exotiny._0022_[2] ),
    .S(net984),
    .X(_01299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07827_ (.A0(net2307),
    .A1(\i_exotiny._0022_[3] ),
    .S(net984),
    .X(_01300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07828_ (.A0(net3119),
    .A1(net2134),
    .S(net987),
    .X(_01301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07829_ (.A0(net3124),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[5] ),
    .S(net986),
    .X(_01302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07830_ (.A0(net3048),
    .A1(net2162),
    .S(net984),
    .X(_01303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07831_ (.A0(net3137),
    .A1(net2307),
    .S(net983),
    .X(_01304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07832_ (.A0(net2808),
    .A1(net3119),
    .S(net986),
    .X(_01305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07833_ (.A0(net3333),
    .A1(net3124),
    .S(net986),
    .X(_01306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07834_ (.A0(net2142),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[10] ),
    .S(net984),
    .X(_01307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07835_ (.A0(net3222),
    .A1(net3137),
    .S(net983),
    .X(_01308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07836_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[16] ),
    .A1(net2808),
    .S(net986),
    .X(_01309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07837_ (.A0(net3254),
    .A1(net3333),
    .S(net986),
    .X(_01310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07838_ (.A0(net2922),
    .A1(net2142),
    .S(net984),
    .X(_01311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07839_ (.A0(net3446),
    .A1(net3222),
    .S(net983),
    .X(_01312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07840_ (.A0(net2469),
    .A1(net3259),
    .S(net986),
    .X(_01313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07841_ (.A0(net2347),
    .A1(net3254),
    .S(net986),
    .X(_01314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07842_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[22] ),
    .A1(net2922),
    .S(net984),
    .X(_01315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07843_ (.A0(net3420),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[19] ),
    .S(net983),
    .X(_01316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07844_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[24] ),
    .A1(net2469),
    .S(net986),
    .X(_01317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07845_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[25] ),
    .A1(net2347),
    .S(net985),
    .X(_01318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07846_ (.A0(net3252),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[22] ),
    .S(net985),
    .X(_01319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07847_ (.A0(net2536),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[23] ),
    .S(net983),
    .X(_01320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07848_ (.A0(net2471),
    .A1(net3134),
    .S(net987),
    .X(_01321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07849_ (.A0(net2910),
    .A1(net3273),
    .S(net983),
    .X(_01322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07850_ (.A0(net2121),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[26] ),
    .S(net984),
    .X(_01323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07851_ (.A0(net2267),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[27] ),
    .S(net983),
    .X(_01324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07852_ (.A0(\i_exotiny._0022_[0] ),
    .A1(net889),
    .S(_03222_),
    .X(_03224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07853_ (.A0(_03224_),
    .A1(net2471),
    .S(net985),
    .X(_01325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07854_ (.A0(\i_exotiny._0022_[1] ),
    .A1(net882),
    .S(_03222_),
    .X(_03225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07855_ (.A0(_03225_),
    .A1(net2910),
    .S(net985),
    .X(_01326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07856_ (.A0(net2273),
    .A1(net879),
    .S(_03222_),
    .X(_03226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07857_ (.A0(_03226_),
    .A1(net2121),
    .S(net984),
    .X(_01327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07858_ (.A0(net2592),
    .A1(net875),
    .S(_03222_),
    .X(_03227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07859_ (.A0(_03227_),
    .A1(net2267),
    .S(net983),
    .X(_01328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07860_ (.A(_02477_),
    .B(_02492_),
    .Y(_03228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _07861_ (.A2(_03228_),
    .A1(net1142),
    .B1(net1163),
    .X(_03229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07862_ (.A0(\i_exotiny._0021_[0] ),
    .A1(net2069),
    .S(net982),
    .X(_01329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07863_ (.A0(\i_exotiny._0021_[1] ),
    .A1(net2371),
    .S(net980),
    .X(_01330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07864_ (.A0(\i_exotiny._0021_[2] ),
    .A1(net2451),
    .S(net981),
    .X(_01331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07865_ (.A0(net2804),
    .A1(net3140),
    .S(net981),
    .X(_01332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07866_ (.A0(net2069),
    .A1(net2684),
    .S(net982),
    .X(_01333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07867_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[5] ),
    .A1(net2365),
    .S(net978),
    .X(_01334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07868_ (.A0(net2451),
    .A1(net3268),
    .S(net981),
    .X(_01335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07869_ (.A0(net3140),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[11] ),
    .S(net981),
    .X(_01336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07870_ (.A0(net2684),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[12] ),
    .S(net979),
    .X(_01337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07871_ (.A0(net2365),
    .A1(net2690),
    .S(net978),
    .X(_01338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07872_ (.A0(net3268),
    .A1(net3445),
    .S(net981),
    .X(_01339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07873_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[11] ),
    .A1(net2188),
    .S(net980),
    .X(_01340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07874_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[12] ),
    .A1(net3473),
    .S(net979),
    .X(_01341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07875_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[13] ),
    .A1(net2211),
    .S(net978),
    .X(_01342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07876_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[14] ),
    .A1(net3250),
    .S(net981),
    .X(_01343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07877_ (.A0(net2188),
    .A1(net2558),
    .S(net980),
    .X(_01344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07878_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[16] ),
    .A1(net2327),
    .S(net979),
    .X(_01345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07879_ (.A0(net2211),
    .A1(net2981),
    .S(net978),
    .X(_01346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07880_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[18] ),
    .A1(net2259),
    .S(net982),
    .X(_01347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07881_ (.A0(net2558),
    .A1(net2938),
    .S(net980),
    .X(_01348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07882_ (.A0(net2327),
    .A1(net2412),
    .S(net979),
    .X(_01349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07883_ (.A0(net2981),
    .A1(net2810),
    .S(net978),
    .X(_01350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07884_ (.A0(net2259),
    .A1(net3150),
    .S(net982),
    .X(_01351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07885_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[23] ),
    .A1(net2190),
    .S(_03229_),
    .X(_01352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07886_ (.A0(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[24] ),
    .A1(net2253),
    .S(net979),
    .X(_01353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07887_ (.A0(net2810),
    .A1(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[29] ),
    .S(net978),
    .X(_01354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07888_ (.A0(net3150),
    .A1(net3066),
    .S(net981),
    .X(_01355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07889_ (.A0(net2190),
    .A1(net2779),
    .S(net980),
    .X(_01356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07890_ (.A0(net2534),
    .A1(net886),
    .S(_03228_),
    .X(_03230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07891_ (.A0(net2253),
    .A1(_03230_),
    .S(net978),
    .X(_01357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07892_ (.A0(\i_exotiny._0021_[1] ),
    .A1(net881),
    .S(_03228_),
    .X(_03231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07893_ (.A0(net3097),
    .A1(_03231_),
    .S(net978),
    .X(_01358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07894_ (.A0(\i_exotiny._0021_[2] ),
    .A1(net876),
    .S(_03228_),
    .X(_03232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07895_ (.A0(net3066),
    .A1(_03232_),
    .S(net981),
    .X(_01359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07896_ (.A0(net2804),
    .A1(net872),
    .S(_03228_),
    .X(_03233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _07897_ (.A0(net2779),
    .A1(_03233_),
    .S(net980),
    .X(_01360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _07898_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1),
    .Q(\i_exotiny.i_rstctl.sys_res_n ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _07899_ (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00001_),
    .Q(\i_exotiny._1312_ ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _07900_ (.RESET_B(net46),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00002_),
    .Q(\i_exotiny._1306_ ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _07901_ (.RESET_B(net47),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00003_),
    .Q(\i_exotiny._1309_ ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _07902_ (.RESET_B(net48),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00000_),
    .Q(\i_exotiny._1429_ ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _07903_ (.RESET_B(net50),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00004_),
    .Q(\i_exotiny._1308_ ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _07904_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3696),
    .Q(\i_exotiny._1311_ ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _07905_ (.RESET_B(net1176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3568),
    .Q(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.genblk7.g_value.r_value [0]),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _07906_ (.RESET_B(\i_exotiny._0000_ ),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1105),
    .Q(\i_exotiny.i_wdg_top.fsm_inst.sw_trg_s1wto ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _07907_ (.RESET_B(net1176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3512),
    .Q(_00014_),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _07908_ (.RESET_B(net1175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1127),
    .Q(\i_exotiny._3871_ ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _07909_ (.RESET_B(net739),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1979),
    .Q(\i_exotiny._1924_[2] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _07910_ (.RESET_B(net738),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1904),
    .Q(\i_exotiny._1924_[3] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _07911_ (.RESET_B(net737),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1908),
    .Q(\i_exotiny._1924_[4] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _07912_ (.RESET_B(net736),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2051),
    .Q(\i_exotiny._1924_[5] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _07913_ (.RESET_B(net735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1988),
    .Q(\i_exotiny._1924_[6] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _07914_ (.RESET_B(net734),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1896),
    .Q(\i_exotiny._1924_[7] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _07915_ (.RESET_B(net733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1942),
    .Q(\i_exotiny._1924_[8] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _07916_ (.RESET_B(net732),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1944),
    .Q(\i_exotiny._1924_[9] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _07917_ (.RESET_B(net731),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2007),
    .Q(\i_exotiny._1924_[10] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _07918_ (.RESET_B(net730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1910),
    .Q(\i_exotiny._1924_[11] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _07919_ (.RESET_B(net729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1923),
    .Q(\i_exotiny._1924_[12] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _07920_ (.RESET_B(net728),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1954),
    .Q(\i_exotiny._1924_[13] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _07921_ (.RESET_B(net727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1940),
    .Q(\i_exotiny._1924_[14] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _07922_ (.RESET_B(net726),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1964),
    .Q(\i_exotiny._1924_[15] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _07923_ (.RESET_B(net725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2005),
    .Q(\i_exotiny._1924_[16] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _07924_ (.RESET_B(net724),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2032),
    .Q(\i_exotiny._1924_[17] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _07925_ (.RESET_B(net723),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1902),
    .Q(\i_exotiny._1924_[18] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _07926_ (.RESET_B(net722),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1948),
    .Q(\i_exotiny._1924_[19] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _07927_ (.RESET_B(net721),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1958),
    .Q(\i_exotiny._1924_[20] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _07928_ (.RESET_B(net720),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1917),
    .Q(\i_exotiny._1924_[21] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _07929_ (.RESET_B(net719),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1927),
    .Q(\i_exotiny._1924_[22] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _07930_ (.RESET_B(net718),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2047),
    .Q(\i_exotiny._1924_[23] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _07931_ (.RESET_B(net717),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2529),
    .Q(\i_exotiny._1924_[24] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _07932_ (.RESET_B(net716),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1921),
    .Q(\i_exotiny._1924_[25] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _07933_ (.RESET_B(net715),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1983),
    .Q(\i_exotiny._1924_[26] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _07934_ (.RESET_B(net714),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1925),
    .Q(\i_exotiny._1924_[27] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _07935_ (.RESET_B(net713),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1919),
    .Q(\i_exotiny._1924_[28] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _07936_ (.RESET_B(net712),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1900),
    .Q(\i_exotiny._1924_[29] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _07937_ (.RESET_B(net711),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1999),
    .Q(\i_exotiny._1924_[30] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _07938_ (.RESET_B(net710),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1960),
    .Q(\i_exotiny._1924_[31] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _07939_ (.RESET_B(net709),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1929),
    .Q(\i_exotiny.i_wb_spi.spi_sdo_o ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _07940_ (.RESET_B(net1175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2034),
    .Q(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.genblk7.g_value.r_value [0]),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _07941_ (.RESET_B(net85),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00006_),
    .Q(\i_exotiny._1793_ ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _07942_ (.RESET_B(net86),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3522),
    .Q(\i_exotiny._1715_ ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _07943_ (.RESET_B(net87),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00008_),
    .Q(\i_exotiny._1737_ ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _07944_ (.RESET_B(net88),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3755),
    .Q(\i_exotiny._1660_ ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _07945_ (.RESET_B(net89),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3653),
    .Q(\i_exotiny._1757_ ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _07946_ (.RESET_B(net90),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00011_),
    .Q(\i_exotiny._1711_ ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _07947_ (.RESET_B(net94),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00012_),
    .Q(\i_exotiny._1725_ ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _07948_ (.RESET_B(net708),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00013_),
    .Q(\i_exotiny._1623_ ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _07949_ (.RESET_B(net707),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1973),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[4] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _07950_ (.RESET_B(net706),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3704),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[5] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _07951_ (.RESET_B(net95),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1932),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[6] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _07952_ (.RESET_B(net1179),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3782),
    .Q(\i_exotiny.i_wdg_top.do_cnt ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _07953_ (.RESET_B(net1179),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1833),
    .Q(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_hw_set [0]),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _07954_ (.RESET_B(net1179),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2055_[2] ),
    .Q(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set [0]),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _07955_ (.RESET_B(net705),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00062_),
    .Q(\i_exotiny._1956_ ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _07956_ (.RESET_B(net703),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00063_),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[1] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _07957_ (.RESET_B(net700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3401),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[2] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _07958_ (.RESET_B(net698),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1993),
    .Q(\i_exotiny.i_wb_spi.cnt_hbit_r[3] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _07959_ (.RESET_B(net1176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3736),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[0] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _07960_ (.RESET_B(net1175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3554),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[1] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _07961_ (.RESET_B(net1176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3667),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[2] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _07962_ (.RESET_B(net1176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3529),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[3] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _07963_ (.RESET_B(net1175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3786),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[4] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _07964_ (.RESET_B(net1175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3797),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[5] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _07965_ (.RESET_B(net1177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3753),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[6] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _07966_ (.RESET_B(net1178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3716),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[7] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _07967_ (.RESET_B(net1178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3710),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[8] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _07968_ (.RESET_B(net1177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3793),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[9] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _07969_ (.RESET_B(net1175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1889),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[10] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _07970_ (.RESET_B(net1177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1871),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[11] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _07971_ (.RESET_B(net1177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1876),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[12] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _07972_ (.RESET_B(net1178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1874),
    .Q(\i_exotiny.i_wdg_top.o_wb_dat[13] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _07973_ (.RESET_B(net114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1611_[1] ),
    .Q(\i_exotiny._0369_[25] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _07974_ (.RESET_B(net115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1611_[2] ),
    .Q(\i_exotiny._0369_[26] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _07975_ (.RESET_B(net116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1611_[3] ),
    .Q(\i_exotiny._0369_[27] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _07976_ (.RESET_B(net117),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3595),
    .Q(\i_exotiny._0369_[29] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _07977_ (.RESET_B(net118),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1611_[6] ),
    .Q(\i_exotiny._0369_[30] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _07978_ (.RESET_B(net119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3585),
    .Q(\i_exotiny._1840_[11] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _07979_ (.RESET_B(net120),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3602),
    .Q(\i_exotiny._0369_[17] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _07980_ (.RESET_B(net121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3458),
    .Q(\i_exotiny._0369_[18] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _07981_ (.RESET_B(net122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3388),
    .Q(\i_exotiny._0369_[19] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_2 _07982_ (.RESET_B(net123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3676),
    .Q(\i_exotiny._0369_[21] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_2 _07983_ (.RESET_B(net124),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3738),
    .Q(\i_exotiny._0369_[22] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_2 _07984_ (.RESET_B(net125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3506),
    .Q(\i_exotiny._0369_[23] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _07985_ (.RESET_B(net126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2126),
    .Q(\i_exotiny._0369_[9] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_2 _07986_ (.RESET_B(net127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3308),
    .Q(\i_exotiny._0369_[10] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_2 _07987_ (.RESET_B(net128),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2062),
    .Q(\i_exotiny._0369_[11] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_2 _07988_ (.RESET_B(net129),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2998),
    .Q(\i_exotiny._0369_[13] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_2 _07989_ (.RESET_B(net130),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3444),
    .Q(\i_exotiny._0369_[14] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_2 _07990_ (.RESET_B(net131),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1611_[23] ),
    .Q(\i_exotiny._0369_[15] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _07991_ (.RESET_B(net132),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3750),
    .Q(\i_exotiny._0369_[1] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _07992_ (.RESET_B(net133),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1611_[26] ),
    .Q(\i_exotiny._0369_[2] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_2 _07993_ (.RESET_B(net134),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3597),
    .Q(\i_exotiny._0369_[3] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _07994_ (.RESET_B(net135),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2736),
    .Q(\i_exotiny._0369_[5] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _07995_ (.RESET_B(net136),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3799),
    .Q(\i_exotiny._0369_[6] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _07996_ (.RESET_B(net137),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1611_[31] ),
    .Q(\i_exotiny._0369_[7] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _07997_ (.RESET_B(\i_exotiny._2032_ ),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net532),
    .Q(\i_exotiny._2044_[1] ),
    .CLK(net1228));
 sg13g2_dfrbpq_2 _07998_ (.RESET_B(\i_exotiny._2032_ ),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2044_[1] ),
    .Q(\i_exotiny.i_wdg_top.cntr_inst.rst_n_sync ),
    .CLK(net1228));
 sg13g2_dfrbpq_2 _07999_ (.RESET_B(net696),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2485),
    .Q(\i_exotiny._0018_[0] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _08000_ (.RESET_B(net695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2816),
    .Q(\i_exotiny._0018_[1] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _08001_ (.RESET_B(net694),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00082_),
    .Q(\i_exotiny._0018_[2] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _08002_ (.RESET_B(net693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2215),
    .Q(\i_exotiny._0018_[3] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _08003_ (.RESET_B(net692),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2086),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _08004_ (.RESET_B(net691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2322),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _08005_ (.RESET_B(net690),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00086_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _08006_ (.RESET_B(net689),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00087_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _08007_ (.RESET_B(net688),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00088_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _08008_ (.RESET_B(net687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00089_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _08009_ (.RESET_B(net686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2599),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _08010_ (.RESET_B(net685),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00091_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _08011_ (.RESET_B(net684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2153),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _08012_ (.RESET_B(net682),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00093_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _08013_ (.RESET_B(net681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2248),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _08014_ (.RESET_B(net680),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2502),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _08015_ (.RESET_B(net679),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00096_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _08016_ (.RESET_B(net678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00097_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _08017_ (.RESET_B(net677),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00098_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _08018_ (.RESET_B(net676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2288),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _08019_ (.RESET_B(net675),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00100_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _08020_ (.RESET_B(net674),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2544),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _08021_ (.RESET_B(net673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00102_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _08022_ (.RESET_B(net672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00103_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _08023_ (.RESET_B(net671),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00104_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _08024_ (.RESET_B(net670),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00105_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _08025_ (.RESET_B(net669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00106_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _08026_ (.RESET_B(net668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2092),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _08027_ (.RESET_B(net667),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00108_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _08028_ (.RESET_B(net666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3371),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _08029_ (.RESET_B(net665),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00110_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _08030_ (.RESET_B(net664),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00111_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _08031_ (.RESET_B(net663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2483),
    .Q(\i_exotiny._0019_[0] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _08032_ (.RESET_B(net662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2129),
    .Q(\i_exotiny._0019_[1] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _08033_ (.RESET_B(net661),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2868),
    .Q(\i_exotiny._0019_[2] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _08034_ (.RESET_B(net660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2896),
    .Q(\i_exotiny._0019_[3] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _08035_ (.RESET_B(net659),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00116_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _08036_ (.RESET_B(net658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00117_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _08037_ (.RESET_B(net657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00118_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _08038_ (.RESET_B(net656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00119_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _08039_ (.RESET_B(net655),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2932),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _08040_ (.RESET_B(net654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2553),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _08041_ (.RESET_B(net653),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2818),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _08042_ (.RESET_B(net652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2904),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _08043_ (.RESET_B(net651),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00124_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _08044_ (.RESET_B(net650),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2884),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _08045_ (.RESET_B(net649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2352),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _08046_ (.RESET_B(net648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00127_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _08047_ (.RESET_B(net647),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2358),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _08048_ (.RESET_B(net646),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2490),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _08049_ (.RESET_B(net645),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2124),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _08050_ (.RESET_B(net644),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2434),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _08051_ (.RESET_B(net643),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00132_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _08052_ (.RESET_B(net642),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2165),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _08053_ (.RESET_B(net641),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00134_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _08054_ (.RESET_B(net640),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00135_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _08055_ (.RESET_B(net639),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00136_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _08056_ (.RESET_B(net638),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00137_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _08057_ (.RESET_B(net637),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00138_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _08058_ (.RESET_B(net636),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00139_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _08059_ (.RESET_B(net635),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3121),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _08060_ (.RESET_B(net634),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2445),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _08061_ (.RESET_B(net633),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2510),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _08062_ (.RESET_B(net632),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2431),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _08063_ (.RESET_B(net631),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2676),
    .Q(\i_exotiny._0020_[0] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_2 _08064_ (.RESET_B(net630),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3030),
    .Q(\i_exotiny._0020_[1] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_2 _08065_ (.RESET_B(net629),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2169),
    .Q(\i_exotiny._0020_[2] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _08066_ (.RESET_B(net628),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3082),
    .Q(\i_exotiny._0020_[3] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _08067_ (.RESET_B(net627),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2320),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _08068_ (.RESET_B(net626),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2419),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _08069_ (.RESET_B(net625),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00150_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _08070_ (.RESET_B(net624),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00151_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _08071_ (.RESET_B(net623),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00152_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _08072_ (.RESET_B(net622),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00153_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _08073_ (.RESET_B(net621),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2970),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _08074_ (.RESET_B(net620),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2823),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _08075_ (.RESET_B(net619),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2793),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _08076_ (.RESET_B(net618),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2171),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _08077_ (.RESET_B(net617),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00158_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _08078_ (.RESET_B(net616),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00159_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _08079_ (.RESET_B(net615),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3284),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _08080_ (.RESET_B(net614),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00161_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _08081_ (.RESET_B(net613),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2407),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _08082_ (.RESET_B(net612),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00163_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _08083_ (.RESET_B(net611),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2235),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _08084_ (.RESET_B(net610),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2459),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _08085_ (.RESET_B(net609),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00166_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _08086_ (.RESET_B(net608),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2457),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _08087_ (.RESET_B(net607),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00168_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _08088_ (.RESET_B(net606),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00169_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _08089_ (.RESET_B(net605),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00170_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _08090_ (.RESET_B(net604),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00171_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _08091_ (.RESET_B(net603),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2813),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _08092_ (.RESET_B(net602),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2773),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _08093_ (.RESET_B(net601),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2478),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _08094_ (.RESET_B(net600),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2506),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _08095_ (.RESET_B(net599),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3418),
    .Q(\i_exotiny._0013_[0] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_2 _08096_ (.RESET_B(net598),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00177_),
    .Q(\i_exotiny._0013_[1] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_2 _08097_ (.RESET_B(net597),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2208),
    .Q(\i_exotiny._0013_[2] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_2 _08098_ (.RESET_B(net596),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00179_),
    .Q(\i_exotiny._0013_[3] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _08099_ (.RESET_B(net595),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00180_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _08100_ (.RESET_B(net594),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2587),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _08101_ (.RESET_B(net593),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00182_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _08102_ (.RESET_B(net592),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2441),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _08103_ (.RESET_B(net591),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2155),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _08104_ (.RESET_B(net590),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00185_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _08105_ (.RESET_B(net589),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2378),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _08106_ (.RESET_B(net588),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00187_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _08107_ (.RESET_B(net587),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00188_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _08108_ (.RESET_B(net586),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2596),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _08109_ (.RESET_B(net585),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00190_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _08110_ (.RESET_B(net584),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00191_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _08111_ (.RESET_B(net583),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2344),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _08112_ (.RESET_B(net582),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3488),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _08113_ (.RESET_B(net581),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00194_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _08114_ (.RESET_B(net580),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00195_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _08115_ (.RESET_B(net579),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00196_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _08116_ (.RESET_B(net578),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2670),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _08117_ (.RESET_B(net577),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3265),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _08118_ (.RESET_B(net576),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2338),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _08119_ (.RESET_B(net575),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2755),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _08120_ (.RESET_B(net574),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00201_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _08121_ (.RESET_B(net573),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2157),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _08122_ (.RESET_B(net572),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2631),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _08123_ (.RESET_B(net571),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3514),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _08124_ (.RESET_B(net570),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00205_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _08125_ (.RESET_B(net569),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00206_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _08126_ (.RESET_B(net568),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00207_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _08127_ (.RESET_B(net1176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3143),
    .Q(_00015_),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _08128_ (.RESET_B(net1178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1981),
    .Q(_00016_),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _08129_ (.RESET_B(net1177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2332),
    .Q(_00017_),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _08130_ (.RESET_B(net1178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2043),
    .Q(_00018_),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_2 _08131_ (.RESET_B(net1177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3560),
    .Q(_00019_),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _08132_ (.RESET_B(net1175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00213_),
    .Q(_00020_),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _08133_ (.RESET_B(net1177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3544),
    .Q(_00021_),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _08134_ (.RESET_B(net1177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2064),
    .Q(_00022_),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_2 _08135_ (.RESET_B(net1178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2013),
    .Q(_00023_),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_2 _08136_ (.RESET_B(net549),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2638),
    .Q(\i_exotiny._0025_[0] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_2 _08137_ (.RESET_B(net548),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3486),
    .Q(\i_exotiny._0025_[1] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_2 _08138_ (.RESET_B(net547),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00219_),
    .Q(\i_exotiny._0025_[2] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_2 _08139_ (.RESET_B(net546),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2514),
    .Q(\i_exotiny._0025_[3] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _08140_ (.RESET_B(net545),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00221_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _08141_ (.RESET_B(net544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00222_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _08142_ (.RESET_B(net543),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00223_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _08143_ (.RESET_B(net542),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00224_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _08144_ (.RESET_B(net541),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00225_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _08145_ (.RESET_B(net540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2605),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _08146_ (.RESET_B(net539),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00227_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _08147_ (.RESET_B(net531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2612),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _08148_ (.RESET_B(net530),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00229_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _08149_ (.RESET_B(net529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00230_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _08150_ (.RESET_B(net528),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2564),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _08151_ (.RESET_B(net527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3061),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _08152_ (.RESET_B(net526),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2221),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _08153_ (.RESET_B(net525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00234_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _08154_ (.RESET_B(net524),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00235_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _08155_ (.RESET_B(net523),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2019),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _08156_ (.RESET_B(net522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2258),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _08157_ (.RESET_B(net521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2392),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _08158_ (.RESET_B(net520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2700),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _08159_ (.RESET_B(net519),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00240_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _08160_ (.RESET_B(net518),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00241_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _08161_ (.RESET_B(net517),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00242_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _08162_ (.RESET_B(net516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2272),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _08163_ (.RESET_B(net515),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00244_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _08164_ (.RESET_B(net514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2589),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _08165_ (.RESET_B(net513),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2796),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _08166_ (.RESET_B(net512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00247_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _08167_ (.RESET_B(net511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2801),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _08168_ (.RESET_B(net510),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2141),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _08169_ (.RESET_B(net508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00250_),
    .Q(\i_exotiny._0038_[0] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_2 _08170_ (.RESET_B(net507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00251_),
    .Q(\i_exotiny._0038_[1] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_2 _08171_ (.RESET_B(net506),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2256),
    .Q(\i_exotiny._0038_[2] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_2 _08172_ (.RESET_B(net505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2304),
    .Q(\i_exotiny._0038_[3] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _08173_ (.RESET_B(net504),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3350),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _08174_ (.RESET_B(net503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00255_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _08175_ (.RESET_B(net502),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00256_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _08176_ (.RESET_B(net501),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00257_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _08177_ (.RESET_B(net500),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00258_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _08178_ (.RESET_B(net499),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2149),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _08179_ (.RESET_B(net498),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00260_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _08180_ (.RESET_B(net497),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00261_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _08181_ (.RESET_B(net496),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2845),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _08182_ (.RESET_B(net495),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00263_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _08183_ (.RESET_B(net494),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2620),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _08184_ (.RESET_B(net493),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2074),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _08185_ (.RESET_B(net492),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00266_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _08186_ (.RESET_B(net491),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3280),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _08187_ (.RESET_B(net490),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2414),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _08188_ (.RESET_B(net489),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00269_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _08189_ (.RESET_B(net488),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2799),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _08190_ (.RESET_B(net487),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2594),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _08191_ (.RESET_B(net486),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00272_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _08192_ (.RESET_B(net485),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2436),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _08193_ (.RESET_B(net484),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2277),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _08194_ (.RESET_B(net483),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2401),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _08195_ (.RESET_B(net482),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00276_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _08196_ (.RESET_B(net481),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00277_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _08197_ (.RESET_B(net480),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00278_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _08198_ (.RESET_B(net479),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00279_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _08199_ (.RESET_B(net478),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2757),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _08200_ (.RESET_B(net477),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00281_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _08201_ (.RESET_B(net476),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3112),
    .Q(\i_exotiny._0037_[0] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_2 _08202_ (.RESET_B(net475),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2318),
    .Q(\i_exotiny._0037_[1] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_2 _08203_ (.RESET_B(net474),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2962),
    .Q(\i_exotiny._0037_[2] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_2 _08204_ (.RESET_B(net473),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2116),
    .Q(\i_exotiny._0037_[3] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _08205_ (.RESET_B(net472),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00286_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _08206_ (.RESET_B(net471),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00287_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _08207_ (.RESET_B(net470),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00288_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _08208_ (.RESET_B(net469),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00289_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _08209_ (.RESET_B(net468),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2763),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _08210_ (.RESET_B(net467),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00291_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _08211_ (.RESET_B(net466),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2692),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _08212_ (.RESET_B(net465),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2603),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _08213_ (.RESET_B(net464),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3015),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _08214_ (.RESET_B(net463),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00295_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _08215_ (.RESET_B(net462),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3451),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _08216_ (.RESET_B(net461),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00297_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _08217_ (.RESET_B(net460),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00298_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _08218_ (.RESET_B(net459),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00299_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _08219_ (.RESET_B(net458),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2262),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _08220_ (.RESET_B(net457),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00301_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _08221_ (.RESET_B(net456),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00302_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _08222_ (.RESET_B(net455),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00303_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _08223_ (.RESET_B(net454),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00304_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _08224_ (.RESET_B(net453),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2334),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _08225_ (.RESET_B(net452),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2710),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _08226_ (.RESET_B(net451),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2390),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _08227_ (.RESET_B(net450),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00308_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _08228_ (.RESET_B(net449),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00309_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _08229_ (.RESET_B(net448),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3303),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _08230_ (.RESET_B(net447),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2683),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _08231_ (.RESET_B(net446),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2665),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _08232_ (.RESET_B(net445),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00313_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_2 _08233_ (.RESET_B(net444),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3128),
    .Q(\i_exotiny._0028_[0] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_2 _08234_ (.RESET_B(net443),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3394),
    .Q(\i_exotiny._0028_[1] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_2 _08235_ (.RESET_B(net442),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2167),
    .Q(\i_exotiny._0028_[2] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _08236_ (.RESET_B(net441),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3103),
    .Q(\i_exotiny._0028_[3] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _08237_ (.RESET_B(net440),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00318_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _08238_ (.RESET_B(net439),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3278),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _08239_ (.RESET_B(net438),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00320_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _08240_ (.RESET_B(net437),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00321_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _08241_ (.RESET_B(net436),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3192),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _08242_ (.RESET_B(net435),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2219),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _08243_ (.RESET_B(net434),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00324_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _08244_ (.RESET_B(net433),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2740),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _08245_ (.RESET_B(net432),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3246),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _08246_ (.RESET_B(net431),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00327_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _08247_ (.RESET_B(net430),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00328_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _08248_ (.RESET_B(net429),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2264),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _08249_ (.RESET_B(net428),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2110),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _08250_ (.RESET_B(net427),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00331_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _08251_ (.RESET_B(net426),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00332_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _08252_ (.RESET_B(net425),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2239),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _08253_ (.RESET_B(net424),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00334_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _08254_ (.RESET_B(net423),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2227),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _08255_ (.RESET_B(net422),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00336_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _08256_ (.RESET_B(net421),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00337_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _08257_ (.RESET_B(net420),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00338_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _08258_ (.RESET_B(net419),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00339_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _08259_ (.RESET_B(net418),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00340_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _08260_ (.RESET_B(net417),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00341_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _08261_ (.RESET_B(net416),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00342_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _08262_ (.RESET_B(net415),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3024),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _08263_ (.RESET_B(net414),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3162),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _08264_ (.RESET_B(net413),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00345_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _08265_ (.RESET_B(net1175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2088),
    .Q(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.genblk7.g_value.r_value [0]),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _08266_ (.RESET_B(net412),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2147),
    .Q(\i_exotiny._0033_[0] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_2 _08267_ (.RESET_B(net411),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2231),
    .Q(\i_exotiny._0033_[1] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_2 _08268_ (.RESET_B(net410),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00349_),
    .Q(\i_exotiny._0033_[2] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_2 _08269_ (.RESET_B(net409),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00350_),
    .Q(\i_exotiny._0033_[3] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _08270_ (.RESET_B(net408),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00351_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _08271_ (.RESET_B(net407),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00352_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _08272_ (.RESET_B(net406),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00353_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _08273_ (.RESET_B(net405),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3496),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _08274_ (.RESET_B(net404),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00355_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _08275_ (.RESET_B(net403),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00356_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _08276_ (.RESET_B(net402),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2428),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _08277_ (.RESET_B(net401),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3480),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _08278_ (.RESET_B(net400),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00359_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _08279_ (.RESET_B(net399),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00360_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _08280_ (.RESET_B(net398),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00361_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _08281_ (.RESET_B(net397),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3189),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _08282_ (.RESET_B(net396),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00363_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _08283_ (.RESET_B(net395),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00364_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _08284_ (.RESET_B(net394),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2567),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _08285_ (.RESET_B(net393),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2476),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _08286_ (.RESET_B(net392),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2376),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _08287_ (.RESET_B(net391),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2370),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _08288_ (.RESET_B(net390),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00369_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _08289_ (.RESET_B(net389),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00370_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _08290_ (.RESET_B(net388),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2480),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _08291_ (.RESET_B(net387),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2306),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _08292_ (.RESET_B(net386),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00373_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _08293_ (.RESET_B(net385),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00374_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _08294_ (.RESET_B(net384),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3456),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _08295_ (.RESET_B(net383),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00376_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _08296_ (.RESET_B(net382),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2672),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _08297_ (.RESET_B(net381),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3209),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _08298_ (.RESET_B(net380),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2096),
    .Q(\i_exotiny._0031_[0] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_2 _08299_ (.RESET_B(net379),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3516),
    .Q(\i_exotiny._0031_[1] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _08300_ (.RESET_B(net378),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00381_),
    .Q(\i_exotiny._0031_[2] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _08301_ (.RESET_B(net377),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2137),
    .Q(\i_exotiny._0031_[3] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _08302_ (.RESET_B(net376),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00383_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _08303_ (.RESET_B(net375),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2417),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _08304_ (.RESET_B(net374),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3088),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _08305_ (.RESET_B(net373),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00386_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _08306_ (.RESET_B(net372),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2987),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _08307_ (.RESET_B(net371),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00388_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _08308_ (.RESET_B(net370),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00389_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _08309_ (.RESET_B(net369),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00390_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _08310_ (.RESET_B(net368),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00391_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _08311_ (.RESET_B(net367),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00392_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _08312_ (.RESET_B(net366),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3286),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _08313_ (.RESET_B(net365),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00394_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _08314_ (.RESET_B(net364),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2622),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _08315_ (.RESET_B(net363),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00396_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _08316_ (.RESET_B(net362),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2181),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _08317_ (.RESET_B(net361),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00398_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _08318_ (.RESET_B(net360),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2201),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _08319_ (.RESET_B(net359),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2374),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _08320_ (.RESET_B(net358),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00401_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _08321_ (.RESET_B(net357),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00402_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _08322_ (.RESET_B(net356),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00403_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _08323_ (.RESET_B(net355),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00404_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _08324_ (.RESET_B(net354),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00405_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _08325_ (.RESET_B(net353),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00406_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _08326_ (.RESET_B(net352),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00407_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _08327_ (.RESET_B(net351),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3165),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _08328_ (.RESET_B(net350),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00409_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _08329_ (.RESET_B(net349),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2641),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _08330_ (.RESET_B(net348),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3180),
    .Q(\i_exotiny._0016_[0] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _08331_ (.RESET_B(net347),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2120),
    .Q(\i_exotiny._0016_[1] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_2 _08332_ (.RESET_B(net346),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3027),
    .Q(\i_exotiny._0016_[2] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_2 _08333_ (.RESET_B(net345),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00414_),
    .Q(\i_exotiny._0016_[3] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _08334_ (.RESET_B(net344),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2403),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _08335_ (.RESET_B(net343),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00416_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _08336_ (.RESET_B(net342),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00417_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _08337_ (.RESET_B(net341),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00418_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _08338_ (.RESET_B(net340),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00419_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _08339_ (.RESET_B(net339),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00420_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _08340_ (.RESET_B(net338),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2776),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _08341_ (.RESET_B(net337),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2386),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _08342_ (.RESET_B(net336),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2508),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _08343_ (.RESET_B(net335),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00424_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _08344_ (.RESET_B(net334),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00425_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _08345_ (.RESET_B(net333),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3406),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _08346_ (.RESET_B(net332),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00427_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _08347_ (.RESET_B(net331),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00428_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _08348_ (.RESET_B(net330),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00429_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _08349_ (.RESET_B(net329),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2821),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _08350_ (.RESET_B(net328),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00431_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _08351_ (.RESET_B(net327),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2368),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _08352_ (.RESET_B(net326),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3230),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _08353_ (.RESET_B(net325),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00434_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _08354_ (.RESET_B(net324),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00435_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _08355_ (.RESET_B(net323),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00436_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _08356_ (.RESET_B(net322),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3207),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _08357_ (.RESET_B(net321),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2674),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _08358_ (.RESET_B(net320),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2384),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _08359_ (.RESET_B(net319),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2425),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _08360_ (.RESET_B(net318),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00441_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _08361_ (.RESET_B(net317),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00442_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _08362_ (.RESET_B(net316),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00443_),
    .Q(\i_exotiny._0014_[0] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_2 _08363_ (.RESET_B(net315),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2466),
    .Q(\i_exotiny._0014_[1] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_2 _08364_ (.RESET_B(net314),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00445_),
    .Q(\i_exotiny._0014_[2] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_2 _08365_ (.RESET_B(net313),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00446_),
    .Q(\i_exotiny._0014_[3] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _08366_ (.RESET_B(net312),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00447_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _08367_ (.RESET_B(net311),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00448_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _08368_ (.RESET_B(net310),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00449_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _08369_ (.RESET_B(net309),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00450_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _08370_ (.RESET_B(net308),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00451_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _08371_ (.RESET_B(net307),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00452_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _08372_ (.RESET_B(net306),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00453_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _08373_ (.RESET_B(net305),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2827),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _08374_ (.RESET_B(net304),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2326),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _08375_ (.RESET_B(net303),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2651),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _08376_ (.RESET_B(net302),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3258),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _08377_ (.RESET_B(net301),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3267),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _08378_ (.RESET_B(net300),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1977),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _08379_ (.RESET_B(net299),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2114),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _08380_ (.RESET_B(net298),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2950),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _08381_ (.RESET_B(net297),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2001),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _08382_ (.RESET_B(net296),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00463_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _08383_ (.RESET_B(net295),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00464_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _08384_ (.RESET_B(net294),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2017),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _08385_ (.RESET_B(net293),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00466_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _08386_ (.RESET_B(net292),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00467_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _08387_ (.RESET_B(net291),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2731),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _08388_ (.RESET_B(net290),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00469_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _08389_ (.RESET_B(net289),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00470_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _08390_ (.RESET_B(net288),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00471_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _08391_ (.RESET_B(net287),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3148),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _08392_ (.RESET_B(net286),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2354),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _08393_ (.RESET_B(net533),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00474_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_2 _08394_ (.RESET_B(net534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1902_[0] ),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[0] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _08395_ (.RESET_B(net535),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1902_[1] ),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[1] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _08396_ (.RESET_B(net536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1902_[2] ),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[2] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _08397_ (.RESET_B(net537),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3552),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[3] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _08398_ (.RESET_B(net538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3619),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[4] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _08399_ (.RESET_B(net683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3562),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[5] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _08400_ (.RESET_B(net285),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3431),
    .Q(\i_exotiny.i_wb_spi.cnt_presc_r[6] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _08401_ (.RESET_B(net284),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2139),
    .Q(\i_exotiny._0035_[0] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_2 _08402_ (.RESET_B(net283),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00476_),
    .Q(\i_exotiny._0035_[1] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_2 _08403_ (.RESET_B(net282),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00477_),
    .Q(\i_exotiny._0035_[2] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_2 _08404_ (.RESET_B(net281),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3540),
    .Q(\i_exotiny._0035_[3] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _08405_ (.RESET_B(net280),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00479_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _08406_ (.RESET_B(net279),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3262),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _08407_ (.RESET_B(net278),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3374),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _08408_ (.RESET_B(net277),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2270),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _08409_ (.RESET_B(net276),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2930),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _08410_ (.RESET_B(net275),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00484_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _08411_ (.RESET_B(net274),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2284),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _08412_ (.RESET_B(net273),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00486_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _08413_ (.RESET_B(net272),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3433),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _08414_ (.RESET_B(net271),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3355),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _08415_ (.RESET_B(net270),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00489_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _08416_ (.RESET_B(net269),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2852),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _08417_ (.RESET_B(net268),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2494),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _08418_ (.RESET_B(net267),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00492_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _08419_ (.RESET_B(net266),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00493_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _08420_ (.RESET_B(net265),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00494_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _08421_ (.RESET_B(net264),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00495_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _08422_ (.RESET_B(net263),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2474),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _08423_ (.RESET_B(net262),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2197),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _08424_ (.RESET_B(net261),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2516),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _08425_ (.RESET_B(net260),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2996),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _08426_ (.RESET_B(net259),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00500_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _08427_ (.RESET_B(net258),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00501_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _08428_ (.RESET_B(net257),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00502_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _08429_ (.RESET_B(net256),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3325),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _08430_ (.RESET_B(net255),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2577),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _08431_ (.RESET_B(net254),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00505_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _08432_ (.RESET_B(net253),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2523),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _08433_ (.RESET_B(net252),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00507_),
    .Q(\i_exotiny._0369_[24] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _08434_ (.RESET_B(net251),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00508_),
    .Q(\i_exotiny._0369_[28] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _08435_ (.RESET_B(net250),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3765),
    .Q(\i_exotiny._0369_[16] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _08436_ (.RESET_B(net249),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00510_),
    .Q(\i_exotiny._0369_[20] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _08437_ (.RESET_B(net248),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00511_),
    .Q(\i_exotiny._0369_[8] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _08438_ (.RESET_B(net247),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3779),
    .Q(\i_exotiny._0369_[12] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _08439_ (.RESET_B(net246),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3760),
    .Q(\i_exotiny._0369_[0] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _08440_ (.RESET_B(net245),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2015),
    .Q(\i_exotiny._0369_[4] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _08441_ (.RESET_B(net244),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00515_),
    .Q(\i_exotiny._2025_[3] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _08442_ (.RESET_B(net242),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00516_),
    .Q(\i_exotiny._2025_[4] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _08443_ (.RESET_B(net240),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00517_),
    .Q(\i_exotiny._2025_[5] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _08444_ (.RESET_B(net238),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00518_),
    .Q(\i_exotiny._2025_[6] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _08445_ (.RESET_B(net236),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00519_),
    .Q(\i_exotiny.i_wb_qspi_mem.crm_r ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _08446_ (.RESET_B(net234),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00520_),
    .Q(\i_exotiny.i_wb_regs.spi_size_o[0] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _08447_ (.RESET_B(net233),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00521_),
    .Q(\i_exotiny.i_wb_regs.spi_size_o[1] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _08448_ (.RESET_B(net232),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2906),
    .Q(\i_exotiny._0039_[0] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_2 _08449_ (.RESET_B(net231),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00523_),
    .Q(\i_exotiny._0039_[1] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_2 _08450_ (.RESET_B(net230),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00524_),
    .Q(\i_exotiny._0039_[2] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_2 _08451_ (.RESET_B(net229),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3345),
    .Q(\i_exotiny._0039_[3] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _08452_ (.RESET_B(net228),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00526_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _08453_ (.RESET_B(net227),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00527_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _08454_ (.RESET_B(net226),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00528_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _08455_ (.RESET_B(net225),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2058),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _08456_ (.RESET_B(net224),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2610),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _08457_ (.RESET_B(net223),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2233),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _08458_ (.RESET_B(net222),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2551),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _08459_ (.RESET_B(net221),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00533_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _08460_ (.RESET_B(net220),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00534_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _08461_ (.RESET_B(net219),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2382),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _08462_ (.RESET_B(net218),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2649),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _08463_ (.RESET_B(net217),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00537_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _08464_ (.RESET_B(net216),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2738),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _08465_ (.RESET_B(net215),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00539_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _08466_ (.RESET_B(net214),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00540_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _08467_ (.RESET_B(net213),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00541_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _08468_ (.RESET_B(net212),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3069),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _08469_ (.RESET_B(net211),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00543_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _08470_ (.RESET_B(net210),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00544_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _08471_ (.RESET_B(net209),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3116),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _08472_ (.RESET_B(net208),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3152),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _08473_ (.RESET_B(net207),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2250),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _08474_ (.RESET_B(net206),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00548_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _08475_ (.RESET_B(net205),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00549_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _08476_ (.RESET_B(net204),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3329),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _08477_ (.RESET_B(net203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00551_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _08478_ (.RESET_B(net202),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00552_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _08479_ (.RESET_B(net201),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3347),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_2 _08480_ (.RESET_B(net200),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00554_),
    .Q(\i_exotiny._0041_[0] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_2 _08481_ (.RESET_B(net199),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00555_),
    .Q(\i_exotiny._0041_[1] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_2 _08482_ (.RESET_B(net198),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3483),
    .Q(\i_exotiny._0041_[2] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_2 _08483_ (.RESET_B(net197),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2082),
    .Q(\i_exotiny._0041_[3] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _08484_ (.RESET_B(net196),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00558_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _08485_ (.RESET_B(net195),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2984),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _08486_ (.RESET_B(net194),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2531),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _08487_ (.RESET_B(net193),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00561_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _08488_ (.RESET_B(net192),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00562_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _08489_ (.RESET_B(net191),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3020),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _08490_ (.RESET_B(net190),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00564_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _08491_ (.RESET_B(net189),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00565_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _08492_ (.RESET_B(net188),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00566_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _08493_ (.RESET_B(net187),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2877),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _08494_ (.RESET_B(net186),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00568_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _08495_ (.RESET_B(net185),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00569_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _08496_ (.RESET_B(net184),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2449),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _08497_ (.RESET_B(net183),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00571_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _08498_ (.RESET_B(net182),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00572_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _08499_ (.RESET_B(net181),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2941),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _08500_ (.RESET_B(net180),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2229),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _08501_ (.RESET_B(net179),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00575_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _08502_ (.RESET_B(net178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00576_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _08503_ (.RESET_B(net177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00577_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _08504_ (.RESET_B(net176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00578_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _08505_ (.RESET_B(net175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00579_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _08506_ (.RESET_B(net174),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00580_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _08507_ (.RESET_B(net173),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2364),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _08508_ (.RESET_B(net172),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00582_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _08509_ (.RESET_B(net171),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2533),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _08510_ (.RESET_B(net170),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2342),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _08511_ (.RESET_B(net169),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3118),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_2 _08512_ (.RESET_B(net168),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00586_),
    .Q(\i_exotiny._0043_[0] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_2 _08513_ (.RESET_B(net167),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2286),
    .Q(\i_exotiny._0043_[1] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_2 _08514_ (.RESET_B(net166),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3095),
    .Q(\i_exotiny._0043_[2] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_2 _08515_ (.RESET_B(net165),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2275),
    .Q(\i_exotiny._0043_[3] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _08516_ (.RESET_B(net164),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2836),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _08517_ (.RESET_B(net163),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00591_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _08518_ (.RESET_B(net162),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2825),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _08519_ (.RESET_B(net161),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00593_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _08520_ (.RESET_B(net160),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3154),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _08521_ (.RESET_B(net159),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00595_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _08522_ (.RESET_B(net158),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00596_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _08523_ (.RESET_B(net157),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00597_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _08524_ (.RESET_B(net156),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2875),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _08525_ (.RESET_B(net155),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00599_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _08526_ (.RESET_B(net154),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2185),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _08527_ (.RESET_B(net153),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2225),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _08528_ (.RESET_B(net152),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2702),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _08529_ (.RESET_B(net151),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3055),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _08530_ (.RESET_B(net150),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00604_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _08531_ (.RESET_B(net149),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00605_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _08532_ (.RESET_B(net148),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00606_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _08533_ (.RESET_B(net147),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2624),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _08534_ (.RESET_B(net146),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00608_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _08535_ (.RESET_B(net145),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00609_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _08536_ (.RESET_B(net144),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2618),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _08537_ (.RESET_B(net143),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2151),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _08538_ (.RESET_B(net142),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2966),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _08539_ (.RESET_B(net141),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00613_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _08540_ (.RESET_B(net140),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00614_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _08541_ (.RESET_B(net139),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00615_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _08542_ (.RESET_B(net138),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3240),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _08543_ (.RESET_B(net113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2492),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _08544_ (.RESET_B(net112),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3592),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _08545_ (.RESET_B(net111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3758),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _08546_ (.RESET_B(net110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00620_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _08547_ (.RESET_B(net109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00621_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_2 _08548_ (.RESET_B(net108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00622_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _08549_ (.RESET_B(net107),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00623_),
    .Q(\i_exotiny._0077_[0] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _08550_ (.RESET_B(net106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00624_),
    .Q(\i_exotiny._0077_[1] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_2 _08551_ (.RESET_B(net105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00625_),
    .Q(\i_exotiny._0077_[2] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _08552_ (.RESET_B(net104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00626_),
    .Q(\i_exotiny._0077_[3] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _08553_ (.RESET_B(net702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00627_),
    .Q(\i_exotiny._0077_[4] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _08554_ (.RESET_B(net103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1207_ ),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _08555_ (.RESET_B(net102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3494),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[0].i_hadd.a_i ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _08556_ (.RESET_B(net100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3604),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3[1].i_hadd.a_i ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _08557_ (.RESET_B(net98),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3408),
    .Q(\i_exotiny._0314_[2] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _08558_ (.RESET_B(net96),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00631_),
    .Q(\i_exotiny._0314_[3] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _08559_ (.RESET_B(net92),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3477),
    .Q(\i_exotiny._0314_[4] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_2 _08560_ (.RESET_B(net84),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3383),
    .Q(\i_exotiny._0314_[5] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _08561_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00634_),
    .Q(\i_exotiny._0314_[6] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _08562_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3518),
    .Q(\i_exotiny._0314_[7] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _08563_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00636_),
    .Q(\i_exotiny._0314_[8] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _08564_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00637_),
    .Q(\i_exotiny._0314_[9] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _08565_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3463),
    .Q(\i_exotiny._0314_[10] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_2 _08566_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3499),
    .Q(\i_exotiny._0314_[11] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _08567_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3448),
    .Q(\i_exotiny._0314_[12] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _08568_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2865),
    .Q(\i_exotiny._0314_[13] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _08569_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3403),
    .Q(\i_exotiny._0314_[14] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _08570_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3244),
    .Q(\i_exotiny._0314_[15] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _08571_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3359),
    .Q(\i_exotiny._0314_[16] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _08572_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00645_),
    .Q(\i_exotiny._0314_[17] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _08573_ (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00646_),
    .Q(\i_exotiny._0314_[18] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _08574_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3156),
    .Q(\i_exotiny._0314_[19] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _08575_ (.RESET_B(net54),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2039),
    .Q(\i_exotiny._0314_[20] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _08576_ (.RESET_B(net52),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2009),
    .Q(\i_exotiny._0314_[21] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _08577_ (.RESET_B(net49),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1966),
    .Q(\i_exotiny._0314_[22] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _08578_ (.RESET_B(net1826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1975),
    .Q(\i_exotiny._0314_[23] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _08579_ (.RESET_B(net1824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00652_),
    .Q(\i_exotiny._0314_[24] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _08580_ (.RESET_B(net1822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00653_),
    .Q(\i_exotiny._0314_[25] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _08581_ (.RESET_B(net1820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00654_),
    .Q(\i_exotiny._0314_[26] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _08582_ (.RESET_B(net1818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00655_),
    .Q(\i_exotiny._0314_[27] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _08583_ (.RESET_B(net1816),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2447),
    .Q(\i_exotiny._0314_[28] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _08584_ (.RESET_B(net1814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2003),
    .Q(\i_exotiny._0314_[29] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _08585_ (.RESET_B(net1812),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3731),
    .Q(\i_exotiny._0314_[30] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _08586_ (.RESET_B(net740),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00659_),
    .Q(\i_exotiny._0314_[31] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _08587_ (.RESET_B(net1810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1265_ ),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_hlt_pc_ccx ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _08588_ (.RESET_B(net1808),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3633),
    .Q(\i_exotiny._6090_[0] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _08589_ (.RESET_B(net1807),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00661_),
    .Q(\i_exotiny._6090_[1] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _08590_ (.RESET_B(net1806),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3720),
    .Q(\i_exotiny._6090_[2] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _08591_ (.RESET_B(net1805),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00663_),
    .Q(\i_exotiny._6090_[3] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _08592_ (.RESET_B(net1804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00664_),
    .Q(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data [0]),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _08593_ (.RESET_B(net1803),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00665_),
    .Q(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data [0]),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _08594_ (.RESET_B(net1802),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00666_),
    .Q(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data [0]),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _08595_ (.RESET_B(net1801),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00667_),
    .Q(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data [0]),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _08596_ (.RESET_B(net1800),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3809),
    .Q(\i_exotiny._1612_[0] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _08597_ (.RESET_B(net1799),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00669_),
    .Q(\i_exotiny._1612_[1] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _08598_ (.RESET_B(net1798),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00670_),
    .Q(\i_exotiny._1612_[2] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _08599_ (.RESET_B(net1797),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00671_),
    .Q(\i_exotiny._1612_[3] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _08600_ (.RESET_B(net1796),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00672_),
    .Q(\i_exotiny._1615_[0] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _08601_ (.RESET_B(net1795),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00673_),
    .Q(\i_exotiny._1615_[1] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _08602_ (.RESET_B(net1794),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00674_),
    .Q(\i_exotiny._1615_[2] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _08603_ (.RESET_B(net1793),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00675_),
    .Q(\i_exotiny._1615_[3] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _08604_ (.RESET_B(net1792),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00676_),
    .Q(\i_exotiny._1614_[0] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _08605_ (.RESET_B(net1791),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00677_),
    .Q(\i_exotiny._1614_[1] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _08606_ (.RESET_B(net1790),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3631),
    .Q(\i_exotiny._1614_[2] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _08607_ (.RESET_B(net1789),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00679_),
    .Q(\i_exotiny._1614_[3] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _08608_ (.RESET_B(net1788),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3718),
    .Q(\i_exotiny._1617_[0] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _08609_ (.RESET_B(net1787),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00681_),
    .Q(\i_exotiny._1617_[1] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _08610_ (.RESET_B(net1786),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3564),
    .Q(\i_exotiny._1617_[2] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _08611_ (.RESET_B(net1785),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00683_),
    .Q(\i_exotiny._1617_[3] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _08612_ (.RESET_B(net1784),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3502),
    .Q(\i_exotiny._1616_[0] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _08613_ (.RESET_B(net1783),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3573),
    .Q(\i_exotiny._1616_[1] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _08614_ (.RESET_B(net1782),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3615),
    .Q(\i_exotiny._1616_[2] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _08615_ (.RESET_B(net1781),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3621),
    .Q(\i_exotiny._1616_[3] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_2 _08616_ (.RESET_B(net1780),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3669),
    .Q(\i_exotiny._1619_[0] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _08617_ (.RESET_B(net1779),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00689_),
    .Q(\i_exotiny._1619_[1] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _08618_ (.RESET_B(net1778),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3673),
    .Q(\i_exotiny._1619_[2] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _08619_ (.RESET_B(net1777),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3748),
    .Q(\i_exotiny._1619_[3] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _08620_ (.RESET_B(net1776),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00692_),
    .Q(\i_exotiny._1618_[0] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _08621_ (.RESET_B(net1775),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00693_),
    .Q(\i_exotiny._1618_[1] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _08622_ (.RESET_B(net1774),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00694_),
    .Q(\i_exotiny._1618_[2] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _08623_ (.RESET_B(net1773),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00695_),
    .Q(\i_exotiny._1618_[3] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _08624_ (.RESET_B(net1772),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3467),
    .Q(\i_exotiny._1586_ ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _08625_ (.RESET_B(net1770),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00697_),
    .Q(\i_exotiny.i_rstctl.wdg_res_n ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _08626_ (.RESET_B(net741),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2572),
    .Q(\i_exotiny.core_res_en_n ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _08627_ (.RESET_B(net742),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3524),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _08628_ (.RESET_B(net743),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3679),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _08629_ (.RESET_B(net774),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1986),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[2] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _08630_ (.RESET_B(net1768),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1489_[3] ),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[3] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _08631_ (.RESET_B(net1766),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2636),
    .Q(\i_exotiny._0029_[0] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_2 _08632_ (.RESET_B(net1765),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2525),
    .Q(\i_exotiny._0029_[1] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_2 _08633_ (.RESET_B(net1764),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2409),
    .Q(\i_exotiny._0029_[2] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_2 _08634_ (.RESET_B(net1763),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00702_),
    .Q(\i_exotiny._0029_[3] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _08635_ (.RESET_B(net1762),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00703_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _08636_ (.RESET_B(net1761),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00704_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _08637_ (.RESET_B(net1760),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00705_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _08638_ (.RESET_B(net1759),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00706_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _08639_ (.RESET_B(net1758),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2689),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _08640_ (.RESET_B(net1757),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2857),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _08641_ (.RESET_B(net1756),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2784),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _08642_ (.RESET_B(net1755),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2849),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _08643_ (.RESET_B(net1754),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3381),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _08644_ (.RESET_B(net1753),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2266),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _08645_ (.RESET_B(net1752),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3300),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _08646_ (.RESET_B(net1751),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3042),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _08647_ (.RESET_B(net1750),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3033),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _08648_ (.RESET_B(net1749),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00716_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _08649_ (.RESET_B(net1748),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2279),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _08650_ (.RESET_B(net1747),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2316),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _08651_ (.RESET_B(net1746),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2193),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _08652_ (.RESET_B(net1745),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00720_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _08653_ (.RESET_B(net1744),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00721_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _08654_ (.RESET_B(net1743),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00722_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _08655_ (.RESET_B(net1742),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00723_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _08656_ (.RESET_B(net1741),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00724_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _08657_ (.RESET_B(net1740),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2928),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _08658_ (.RESET_B(net1739),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00726_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _08659_ (.RESET_B(net1738),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00727_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _08660_ (.RESET_B(net1737),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00728_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _08661_ (.RESET_B(net1736),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00729_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _08662_ (.RESET_B(net775),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00730_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_2 _08663_ (.RESET_B(net1203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[0] ),
    .Q(\i_exotiny._2034_[0] ),
    .CLK(net1228));
 sg13g2_dfrbpq_2 _08664_ (.RESET_B(net1203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[1] ),
    .Q(\i_exotiny._2034_[1] ),
    .CLK(net1228));
 sg13g2_dfrbpq_2 _08665_ (.RESET_B(net1203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[2] ),
    .Q(\i_exotiny._2034_[2] ),
    .CLK(net1228));
 sg13g2_dfrbpq_2 _08666_ (.RESET_B(net1203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[3] ),
    .Q(\i_exotiny._2034_[3] ),
    .CLK(net1228));
 sg13g2_dfrbpq_2 _08667_ (.RESET_B(\i_exotiny.i_wdg_top.cntr_inst.rst_n_sync ),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[4] ),
    .Q(\i_exotiny._2034_[4] ),
    .CLK(net1229));
 sg13g2_dfrbpq_2 _08668_ (.RESET_B(\i_exotiny.i_wdg_top.cntr_inst.rst_n_sync ),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[5] ),
    .Q(\i_exotiny._2034_[5] ),
    .CLK(net1229));
 sg13g2_dfrbpq_2 _08669_ (.RESET_B(net1203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[6] ),
    .Q(\i_exotiny._2034_[6] ),
    .CLK(net1229));
 sg13g2_dfrbpq_2 _08670_ (.RESET_B(net1203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[7] ),
    .Q(\i_exotiny._2034_[7] ),
    .CLK(net1229));
 sg13g2_dfrbpq_2 _08671_ (.RESET_B(net1203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[8] ),
    .Q(\i_exotiny._2034_[8] ),
    .CLK(net1229));
 sg13g2_dfrbpq_2 _08672_ (.RESET_B(net1203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._2043_[9] ),
    .Q(\i_exotiny._2034_[9] ),
    .CLK(net1229));
 sg13g2_dfrbpq_2 _08673_ (.RESET_B(net1735),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00731_),
    .Q(\i_exotiny._0034_[0] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_2 _08674_ (.RESET_B(net1734),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2678),
    .Q(\i_exotiny._0034_[1] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_2 _08675_ (.RESET_B(net1733),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2244),
    .Q(\i_exotiny._0034_[2] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_2 _08676_ (.RESET_B(net1732),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00734_),
    .Q(\i_exotiny._0034_[3] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _08677_ (.RESET_B(net1731),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3310),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _08678_ (.RESET_B(net1730),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00736_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _08679_ (.RESET_B(net1729),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00737_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _08680_ (.RESET_B(net1728),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3248),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _08681_ (.RESET_B(net1727),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3100),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _08682_ (.RESET_B(net1726),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00740_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _08683_ (.RESET_B(net1725),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3217),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _08684_ (.RESET_B(net1724),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3289),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _08685_ (.RESET_B(net1723),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2723),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _08686_ (.RESET_B(net1722),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2989),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _08687_ (.RESET_B(net1721),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2330),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _08688_ (.RESET_B(net1720),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2281),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _08689_ (.RESET_B(net1719),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00747_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _08690_ (.RESET_B(net1718),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1995),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _08691_ (.RESET_B(net1717),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00749_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _08692_ (.RESET_B(net1716),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00750_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _08693_ (.RESET_B(net1715),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2909),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _08694_ (.RESET_B(net1714),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00752_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _08695_ (.RESET_B(net1713),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2771),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _08696_ (.RESET_B(net1712),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2926),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _08697_ (.RESET_B(net1711),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2356),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _08698_ (.RESET_B(net1710),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00756_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _08699_ (.RESET_B(net1709),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2161),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _08700_ (.RESET_B(net1708),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2179),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _08701_ (.RESET_B(net1707),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00759_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _08702_ (.RESET_B(net1706),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00760_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _08703_ (.RESET_B(net1705),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00761_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _08704_ (.RESET_B(net1704),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00762_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_2 _08705_ (.RESET_B(net1703),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2060),
    .Q(\i_exotiny._0032_[0] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_2 _08706_ (.RESET_B(net1702),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00764_),
    .Q(\i_exotiny._0032_[1] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_2 _08707_ (.RESET_B(net1701),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2628),
    .Q(\i_exotiny._0032_[2] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_2 _08708_ (.RESET_B(net1700),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2094),
    .Q(\i_exotiny._0032_[3] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _08709_ (.RESET_B(net1699),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00767_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _08710_ (.RESET_B(net1698),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2090),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _08711_ (.RESET_B(net1697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00769_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _08712_ (.RESET_B(net1696),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00770_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _08713_ (.RESET_B(net1695),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00771_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _08714_ (.RESET_B(net1694),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00772_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _08715_ (.RESET_B(net1693),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3035),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _08716_ (.RESET_B(net1692),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00774_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _08717_ (.RESET_B(net1691),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00775_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _08718_ (.RESET_B(net1690),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2076),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _08719_ (.RESET_B(net1689),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00777_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _08720_ (.RESET_B(net1688),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00778_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _08721_ (.RESET_B(net1687),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2646),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _08722_ (.RESET_B(net1686),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00780_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _08723_ (.RESET_B(net1685),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00781_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _08724_ (.RESET_B(net1684),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2913),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _08725_ (.RESET_B(net1683),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3396),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _08726_ (.RESET_B(net1682),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00784_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _08727_ (.RESET_B(net1681),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2112),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _08728_ (.RESET_B(net1680),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3184),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _08729_ (.RESET_B(net1679),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2084),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _08730_ (.RESET_B(net1678),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00788_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _08731_ (.RESET_B(net1677),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00789_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _08732_ (.RESET_B(net1676),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00790_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _08733_ (.RESET_B(net1675),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00791_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _08734_ (.RESET_B(net1674),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00792_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _08735_ (.RESET_B(net1673),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3078),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _08736_ (.RESET_B(net1672),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00794_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_2 _08737_ (.RESET_B(net1671),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2411),
    .Q(\i_exotiny._0017_[0] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _08738_ (.RESET_B(net1670),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00796_),
    .Q(\i_exotiny._0017_[1] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _08739_ (.RESET_B(net1669),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00797_),
    .Q(\i_exotiny._0017_[2] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_2 _08740_ (.RESET_B(net1668),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00798_),
    .Q(\i_exotiny._0017_[3] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _08741_ (.RESET_B(net1667),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00799_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _08742_ (.RESET_B(net1666),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2294),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _08743_ (.RESET_B(net1665),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2921),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _08744_ (.RESET_B(net1664),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3110),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _08745_ (.RESET_B(net1663),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2549),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _08746_ (.RESET_B(net1662),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1829),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _08747_ (.RESET_B(net1661),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00805_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _08748_ (.RESET_B(net1660),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00806_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _08749_ (.RESET_B(net1659),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2394),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _08750_ (.RESET_B(net1658),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00808_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[13] ),
    .CLK(clknet_5_30__leaf_clk_regs));
 sg13g2_dfrbpq_1 _08751_ (.RESET_B(net1657),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00809_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _08752_ (.RESET_B(net1656),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3200),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _08753_ (.RESET_B(net1655),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00811_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _08754_ (.RESET_B(net1654),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2223),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _08755_ (.RESET_B(net1653),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3046),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _08756_ (.RESET_B(net1652),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3426),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _08757_ (.RESET_B(net1651),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2831),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _08758_ (.RESET_B(net1650),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2574),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _08759_ (.RESET_B(net1649),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3276),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _08760_ (.RESET_B(net1648),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2556),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _08761_ (.RESET_B(net1647),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00819_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _08762_ (.RESET_B(net1646),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2807),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _08763_ (.RESET_B(net1645),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2314),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _08764_ (.RESET_B(net1644),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00822_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _08765_ (.RESET_B(net1643),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3305),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _08766_ (.RESET_B(net1642),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00824_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _08767_ (.RESET_B(net1641),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00825_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _08768_ (.RESET_B(net1640),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00826_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _08769_ (.RESET_B(net1639),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00827_),
    .Q(\i_exotiny._0015_[0] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_2 _08770_ (.RESET_B(net1638),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3369),
    .Q(\i_exotiny._0015_[1] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_2 _08771_ (.RESET_B(net1637),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00829_),
    .Q(\i_exotiny._0015_[2] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_2 _08772_ (.RESET_B(net1636),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2360),
    .Q(\i_exotiny._0015_[3] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _08773_ (.RESET_B(net1635),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3001),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _08774_ (.RESET_B(net1634),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3040),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _08775_ (.RESET_B(net1633),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3074),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _08776_ (.RESET_B(net1632),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00834_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _08777_ (.RESET_B(net1631),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00835_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _08778_ (.RESET_B(net1630),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2145),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _08779_ (.RESET_B(net1629),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3365),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _08780_ (.RESET_B(net1628),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00838_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _08781_ (.RESET_B(net1627),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00839_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _08782_ (.RESET_B(net1626),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00840_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _08783_ (.RESET_B(net1625),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00841_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _08784_ (.RESET_B(net1624),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3331),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _08785_ (.RESET_B(net1623),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2968),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _08786_ (.RESET_B(net1622),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2159),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _08787_ (.RESET_B(net1621),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00845_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _08788_ (.RESET_B(net1620),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2118),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _08789_ (.RESET_B(net1619),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3414),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _08790_ (.RESET_B(net1618),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00848_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _08791_ (.RESET_B(net1617),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00849_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _08792_ (.RESET_B(net1616),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00850_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _08793_ (.RESET_B(net1615),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2695),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _08794_ (.RESET_B(net1614),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00852_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _08795_ (.RESET_B(net1613),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3465),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _08796_ (.RESET_B(net1612),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2217),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _08797_ (.RESET_B(net1611),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00855_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _08798_ (.RESET_B(net1610),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2937),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _08799_ (.RESET_B(net1609),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00857_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _08800_ (.RESET_B(net1608),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00858_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_2 _08801_ (.RESET_B(net1607),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3635),
    .Q(\i_exotiny.i_wb_spi.state_r[0] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _08802_ (.RESET_B(net1606),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00860_),
    .Q(\i_exotiny.i_wb_spi.state_r[1] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _08803_ (.RESET_B(net1605),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00861_),
    .Q(\i_exotiny.i_wb_spi.state_r[2] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _08804_ (.RESET_B(net1604),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00862_),
    .Q(\i_exotiny.i_wb_spi.state_r[3] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _08805_ (.RESET_B(net1603),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00863_),
    .Q(\i_exotiny.i_wb_spi.state_r[4] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _08806_ (.RESET_B(net1602),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00864_),
    .Q(\i_exotiny.i_wb_spi.state_r[5] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _08807_ (.RESET_B(net1601),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00865_),
    .Q(\i_exotiny.i_wb_spi.state_r[6] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _08808_ (.RESET_B(net1600),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00866_),
    .Q(\i_exotiny.i_wb_spi.state_r[7] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _08809_ (.RESET_B(net1599),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00867_),
    .Q(\i_exotiny.i_wb_spi.state_r[8] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _08810_ (.RESET_B(net1598),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00868_),
    .Q(\i_exotiny.i_wb_spi.state_r[9] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _08811_ (.RESET_B(net1597),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00869_),
    .Q(\i_exotiny.i_wb_spi.state_r[10] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _08812_ (.RESET_B(net1596),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00870_),
    .Q(\i_exotiny.i_wb_spi.state_r[11] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _08813_ (.RESET_B(net1595),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1850),
    .Q(\i_exotiny.i_wb_spi.state_r[12] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _08814_ (.RESET_B(net1594),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00872_),
    .Q(\i_exotiny.i_wb_spi.state_r[13] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _08815_ (.RESET_B(net1593),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1836),
    .Q(\i_exotiny.i_wb_spi.state_r[14] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _08816_ (.RESET_B(net1592),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1842),
    .Q(\i_exotiny.i_wb_spi.state_r[15] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _08817_ (.RESET_B(net1591),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00875_),
    .Q(\i_exotiny.i_wb_spi.state_r[16] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _08818_ (.RESET_B(net1590),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1860),
    .Q(\i_exotiny.i_wb_spi.state_r[17] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _08819_ (.RESET_B(net1589),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00877_),
    .Q(\i_exotiny.i_wb_spi.state_r[18] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _08820_ (.RESET_B(net1588),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00878_),
    .Q(\i_exotiny.i_wb_spi.state_r[19] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _08821_ (.RESET_B(net1587),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00879_),
    .Q(\i_exotiny.i_wb_spi.state_r[20] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _08822_ (.RESET_B(net1586),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00880_),
    .Q(\i_exotiny.i_wb_spi.state_r[21] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _08823_ (.RESET_B(net1585),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00881_),
    .Q(\i_exotiny.i_wb_spi.state_r[22] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _08824_ (.RESET_B(net1584),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00882_),
    .Q(\i_exotiny.i_wb_spi.state_r[23] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _08825_ (.RESET_B(net1583),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00883_),
    .Q(\i_exotiny.i_wb_spi.state_r[24] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _08826_ (.RESET_B(net1582),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00884_),
    .Q(\i_exotiny.i_wb_spi.state_r[25] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _08827_ (.RESET_B(net1581),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00885_),
    .Q(\i_exotiny.i_wb_spi.state_r[26] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _08828_ (.RESET_B(net1580),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00886_),
    .Q(\i_exotiny.i_wb_spi.state_r[27] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _08829_ (.RESET_B(net1579),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00887_),
    .Q(\i_exotiny.i_wb_spi.state_r[28] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _08830_ (.RESET_B(net1578),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00888_),
    .Q(\i_exotiny.i_wb_spi.state_r[29] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _08831_ (.RESET_B(net1577),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00889_),
    .Q(\i_exotiny.i_wb_spi.state_r[30] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _08832_ (.RESET_B(net1576),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00890_),
    .Q(\i_exotiny.i_wb_spi.state_r[31] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _08833_ (.RESET_B(net1575),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2175),
    .Q(\i_exotiny._0036_[0] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_2 _08834_ (.RESET_B(net1574),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2205),
    .Q(\i_exotiny._0036_[1] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_2 _08835_ (.RESET_B(net1573),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00893_),
    .Q(\i_exotiny._0036_[2] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_2 _08836_ (.RESET_B(net1572),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2080),
    .Q(\i_exotiny._0036_[3] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _08837_ (.RESET_B(net1569),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00895_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _08838_ (.RESET_B(net1568),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00896_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _08839_ (.RESET_B(net1567),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00897_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _08840_ (.RESET_B(net1566),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00898_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _08841_ (.RESET_B(net1565),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2653),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _08842_ (.RESET_B(net1564),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2829),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _08843_ (.RESET_B(net1563),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2788),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _08844_ (.RESET_B(net1562),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00902_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _08845_ (.RESET_B(net1561),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2324),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _08846_ (.RESET_B(net1560),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2199),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _08847_ (.RESET_B(net1559),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3215),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _08848_ (.RESET_B(net1558),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00906_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _08849_ (.RESET_B(net1557),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00907_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _08850_ (.RESET_B(net1556),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00908_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _08851_ (.RESET_B(net1555),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2053),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _08852_ (.RESET_B(net1554),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00910_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _08853_ (.RESET_B(net1553),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00911_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _08854_ (.RESET_B(net1552),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00912_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _08855_ (.RESET_B(net1551),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00913_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _08856_ (.RESET_B(net1550),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2443),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _08857_ (.RESET_B(net1549),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2712),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _08858_ (.RESET_B(net1548),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00916_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _08859_ (.RESET_B(net1547),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00917_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _08860_ (.RESET_B(net1546),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2957),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _08861_ (.RESET_B(net1545),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3534),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _08862_ (.RESET_B(net1544),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2661),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _08863_ (.RESET_B(net1543),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00921_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _08864_ (.RESET_B(net1542),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3438),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _08865_ (.RESET_B(net1541),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00923_),
    .Q(\i_exotiny.i_wb_regs.spi_auto_cs_o ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _08866_ (.RESET_B(net1540),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2108),
    .Q(\i_exotiny.i_wb_regs.spi_cpol_o ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _08867_ (.RESET_B(net1538),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3774),
    .Q(\i_exotiny.gpo[0] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _08868_ (.RESET_B(net1536),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3743),
    .Q(\i_exotiny.gpo[1] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _08869_ (.RESET_B(net1534),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3746),
    .Q(\i_exotiny.gpo[2] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _08870_ (.RESET_B(net1532),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00928_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[0] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _08871_ (.RESET_B(net1531),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3590),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[1] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _08872_ (.RESET_B(net1530),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3577),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[2] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _08873_ (.RESET_B(net1529),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3575),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[3] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _08874_ (.RESET_B(net1528),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3557),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[4] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _08875_ (.RESET_B(net1527),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00933_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[5] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _08876_ (.RESET_B(net1526),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00934_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[6] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _08877_ (.RESET_B(net1525),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1936),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[7] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _08878_ (.RESET_B(net1524),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1969),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[8] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _08879_ (.RESET_B(net1523),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1934),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[9] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _08880_ (.RESET_B(net1522),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00938_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[10] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _08881_ (.RESET_B(net1521),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00939_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[11] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _08882_ (.RESET_B(net1520),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1898),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[12] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _08883_ (.RESET_B(net1519),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1906),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[13] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _08884_ (.RESET_B(net1518),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1946),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[14] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _08885_ (.RESET_B(net1517),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00943_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[15] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _08886_ (.RESET_B(net1516),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00944_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[16] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _08887_ (.RESET_B(net1515),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1952),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[17] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _08888_ (.RESET_B(net1514),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1938),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[18] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _08889_ (.RESET_B(net1513),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00947_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[19] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _08890_ (.RESET_B(net1512),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3645),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[20] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _08891_ (.RESET_B(net1511),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00949_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[21] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _08892_ (.RESET_B(net1510),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00950_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[22] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _08893_ (.RESET_B(net1509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3588),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[23] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _08894_ (.RESET_B(net1508),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3639),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[24] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _08895_ (.RESET_B(net1507),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3664),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[25] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _08896_ (.RESET_B(net1506),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3660),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[26] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _08897_ (.RESET_B(net1505),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3617),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[27] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _08898_ (.RESET_B(net1504),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00956_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[28] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _08899_ (.RESET_B(net1503),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00957_),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[29] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _08900_ (.RESET_B(net1502),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3583),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[30] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _08901_ (.RESET_B(net1501),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3531),
    .Q(\i_exotiny.i_wb_spi.dat_rx_r[31] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_2 _08902_ (.RESET_B(net1500),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00960_),
    .Q(\i_exotiny._0040_[0] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_2 _08903_ (.RESET_B(net1499),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2890),
    .Q(\i_exotiny._0040_[1] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_2 _08904_ (.RESET_B(net1498),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3084),
    .Q(\i_exotiny._0040_[2] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _08905_ (.RESET_B(net1497),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00963_),
    .Q(\i_exotiny._0040_[3] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _08906_ (.RESET_B(net1496),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3315),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _08907_ (.RESET_B(net1495),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00965_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _08908_ (.RESET_B(net1494),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2362),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _08909_ (.RESET_B(net1493),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2468),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _08910_ (.RESET_B(net1492),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2879),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _08911_ (.RESET_B(net1491),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00969_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _08912_ (.RESET_B(net1490),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00970_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _08913_ (.RESET_B(net1489),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00971_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _08914_ (.RESET_B(net1488),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2312),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _08915_ (.RESET_B(net1487),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00973_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _08916_ (.RESET_B(net1486),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2340),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _08917_ (.RESET_B(net1485),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3353),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _08918_ (.RESET_B(net1484),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2310),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _08919_ (.RESET_B(net1483),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00977_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _08920_ (.RESET_B(net1482),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00978_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _08921_ (.RESET_B(net1481),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2455),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _08922_ (.RESET_B(net1480),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00980_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _08923_ (.RESET_B(net1479),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2714),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _08924_ (.RESET_B(net1478),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00982_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _08925_ (.RESET_B(net1477),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00983_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _08926_ (.RESET_B(net1476),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2760),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _08927_ (.RESET_B(net1475),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00985_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _08928_ (.RESET_B(net1474),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00986_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _08929_ (.RESET_B(net1473),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00987_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _08930_ (.RESET_B(net1472),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3072),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _08931_ (.RESET_B(net1471),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2399),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _08932_ (.RESET_B(net1470),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2615),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _08933_ (.RESET_B(net1469),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00991_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_2 _08934_ (.RESET_B(net1468),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2439),
    .Q(\i_exotiny._0042_[0] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _08935_ (.RESET_B(net1467),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00993_),
    .Q(\i_exotiny._0042_[1] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _08936_ (.RESET_B(net1466),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00994_),
    .Q(\i_exotiny._0042_[2] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _08937_ (.RESET_B(net1465),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2203),
    .Q(\i_exotiny._0042_[3] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _08938_ (.RESET_B(net1464),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00996_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _08939_ (.RESET_B(net1463),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2655),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _08940_ (.RESET_B(net1462),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2585),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _08941_ (.RESET_B(net1461),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00999_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _08942_ (.RESET_B(net1460),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01000_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _08943_ (.RESET_B(net1459),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2068),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _08944_ (.RESET_B(net1458),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01002_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _08945_ (.RESET_B(net1457),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2790),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _08946_ (.RESET_B(net1456),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2716),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _08947_ (.RESET_B(net1455),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01005_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _08948_ (.RESET_B(net1454),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2036),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _08949_ (.RESET_B(net1453),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01007_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _08950_ (.RESET_B(net1452),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2246),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _08951_ (.RESET_B(net1451),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01009_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _08952_ (.RESET_B(net1450),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01010_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _08953_ (.RESET_B(net1449),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2847),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _08954_ (.RESET_B(net1448),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01012_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _08955_ (.RESET_B(net1447),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2104),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _08956_ (.RESET_B(net1446),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01014_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _08957_ (.RESET_B(net1445),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3472),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _08958_ (.RESET_B(net1444),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2663),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _08959_ (.RESET_B(net1443),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01017_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _08960_ (.RESET_B(net1442),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2291),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _08961_ (.RESET_B(net1441),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2496),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _08962_ (.RESET_B(net1440),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3233),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _08963_ (.RESET_B(net1439),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01021_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _08964_ (.RESET_B(net1438),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01022_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _08965_ (.RESET_B(net1437),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01023_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _08966_ (.RESET_B(net1436),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01024_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[2] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _08967_ (.RESET_B(net1435),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3691),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[3] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _08968_ (.RESET_B(net1434),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3769),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[4] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _08969_ (.RESET_B(net1433),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01027_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[5] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _08970_ (.RESET_B(net1432),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3685),
    .Q(\i_exotiny._0590_ ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _08971_ (.RESET_B(net1431),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01029_),
    .Q(\i_exotiny._0542_ ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _08972_ (.RESET_B(net1430),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01030_),
    .Q(\i_exotiny._0601_ ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _08973_ (.RESET_B(net1429),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01031_),
    .Q(\i_exotiny._0571_ ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _08974_ (.RESET_B(net1428),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01032_),
    .Q(\i_exotiny._0550_ ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_2 _08975_ (.RESET_B(net1427),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3740),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_2 _08976_ (.RESET_B(net1426),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01034_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _08977_ (.RESET_B(net1425),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01035_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_2 _08978_ (.RESET_B(net1424),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01036_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _08979_ (.RESET_B(net1423),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01037_),
    .Q(\i_exotiny._1160_[0] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _08980_ (.RESET_B(net1422),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2045),
    .Q(\i_exotiny._1160_[1] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _08981_ (.RESET_B(net1421),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01039_),
    .Q(\i_exotiny._1160_[2] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _08982_ (.RESET_B(net1420),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1950),
    .Q(\i_exotiny._1160_[3] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _08983_ (.RESET_B(net1419),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1990),
    .Q(\i_exotiny._1160_[4] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _08984_ (.RESET_B(net1418),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1997),
    .Q(\i_exotiny._1160_[5] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _08985_ (.RESET_B(net1417),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2027),
    .Q(\i_exotiny._1160_[6] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _08986_ (.RESET_B(net1416),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1956),
    .Q(\i_exotiny._1160_[7] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _08987_ (.RESET_B(net1415),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2023),
    .Q(\i_exotiny._1160_[8] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _08988_ (.RESET_B(net1414),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2066),
    .Q(\i_exotiny._1160_[9] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _08989_ (.RESET_B(net1413),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2102),
    .Q(\i_exotiny._1160_[10] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _08990_ (.RESET_B(net1412),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3527),
    .Q(\i_exotiny._1160_[11] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _08991_ (.RESET_B(net1411),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2078),
    .Q(\i_exotiny._1160_[12] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _08992_ (.RESET_B(net1410),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2011),
    .Q(\i_exotiny._1160_[13] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _08993_ (.RESET_B(net1409),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2041),
    .Q(\i_exotiny._1160_[14] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _08994_ (.RESET_B(net1408),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2021),
    .Q(\i_exotiny._1160_[15] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _08995_ (.RESET_B(net1407),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3542),
    .Q(\i_exotiny._1160_[16] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _08996_ (.RESET_B(net1406),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01054_),
    .Q(\i_exotiny._1160_[17] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _08997_ (.RESET_B(net1405),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3566),
    .Q(\i_exotiny._1160_[18] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _08998_ (.RESET_B(net1404),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01056_),
    .Q(\i_exotiny._1160_[19] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _08999_ (.RESET_B(net1403),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3599),
    .Q(\i_exotiny._1160_[20] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _09000_ (.RESET_B(net1402),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3536),
    .Q(\i_exotiny._1160_[21] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _09001_ (.RESET_B(net1401),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01059_),
    .Q(\i_exotiny._1160_[22] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09002_ (.RESET_B(net1400),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01060_),
    .Q(\i_exotiny._1160_[23] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _09003_ (.RESET_B(net1399),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3385),
    .Q(\i_exotiny._1160_[24] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _09004_ (.RESET_B(net1398),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3361),
    .Q(\i_exotiny._1160_[25] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _09005_ (.RESET_B(net1397),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3416),
    .Q(\i_exotiny._1160_[26] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _09006_ (.RESET_B(net1396),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1912),
    .Q(\i_exotiny._1160_[27] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _09007_ (.RESET_B(net1395),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01065_),
    .Q(\i_exotiny._0079_[0] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _09008_ (.RESET_B(net1394),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01066_),
    .Q(\i_exotiny._0079_[1] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_2 _09009_ (.RESET_B(net1393),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01067_),
    .Q(\i_exotiny._0079_[2] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_2 _09010_ (.RESET_B(net1392),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01068_),
    .Q(\i_exotiny._0079_[3] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _09011_ (.RESET_B(net1391),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3581),
    .Q(\i_exotiny._0079_[4] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_2 _09012_ (.RESET_B(net1390),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01070_),
    .Q(\i_exotiny._0327_[0] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _09013_ (.RESET_B(net1389),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01071_),
    .Q(\i_exotiny._0327_[1] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _09014_ (.RESET_B(net1388),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3823),
    .Q(\i_exotiny._0315_[2] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _09015_ (.RESET_B(net1387),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01073_),
    .Q(\i_exotiny._0315_[3] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _09016_ (.RESET_B(net1386),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01074_),
    .Q(\i_exotiny._0315_[4] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _09017_ (.RESET_B(net1385),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01075_),
    .Q(\i_exotiny._0315_[5] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _09018_ (.RESET_B(net1384),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3538),
    .Q(\i_exotiny._0315_[6] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _09019_ (.RESET_B(net1383),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3693),
    .Q(\i_exotiny._0315_[7] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _09020_ (.RESET_B(net1382),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01078_),
    .Q(\i_exotiny._0315_[8] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _09021_ (.RESET_B(net1381),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01079_),
    .Q(\i_exotiny._0315_[9] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _09022_ (.RESET_B(net1380),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01080_),
    .Q(\i_exotiny._0315_[10] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_2 _09023_ (.RESET_B(net1379),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01081_),
    .Q(\i_exotiny._0315_[11] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _09024_ (.RESET_B(net1378),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01082_),
    .Q(\i_exotiny._0315_[12] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _09025_ (.RESET_B(net1377),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3546),
    .Q(\i_exotiny._0315_[13] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _09026_ (.RESET_B(net1376),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3548),
    .Q(\i_exotiny._0315_[14] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09027_ (.RESET_B(net1375),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3613),
    .Q(\i_exotiny._0315_[15] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _09028_ (.RESET_B(net1374),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3662),
    .Q(\i_exotiny._0315_[16] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _09029_ (.RESET_B(net1373),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01087_),
    .Q(\i_exotiny._0315_[17] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _09030_ (.RESET_B(net1372),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3550),
    .Q(\i_exotiny._0315_[18] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09031_ (.RESET_B(net1371),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01089_),
    .Q(\i_exotiny._0315_[19] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _09032_ (.RESET_B(net1370),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2842),
    .Q(\i_exotiny._0315_[20] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _09033_ (.RESET_B(net1369),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01091_),
    .Q(\i_exotiny._0315_[21] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _09034_ (.RESET_B(net1368),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3114),
    .Q(\i_exotiny._0315_[22] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _09035_ (.RESET_B(net1367),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01093_),
    .Q(\i_exotiny._0315_[23] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _09036_ (.RESET_B(net1366),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01094_),
    .Q(\i_exotiny._0315_[24] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _09037_ (.RESET_B(net1365),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3221),
    .Q(\i_exotiny._0315_[25] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _09038_ (.RESET_B(net1364),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01096_),
    .Q(\i_exotiny._0315_[26] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _09039_ (.RESET_B(net1363),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01097_),
    .Q(\i_exotiny._0315_[27] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _09040_ (.RESET_B(net1362),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2100),
    .Q(\i_exotiny._0315_[28] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _09041_ (.RESET_B(net1361),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01099_),
    .Q(\i_exotiny._0315_[29] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _09042_ (.RESET_B(net1360),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01100_),
    .Q(\i_exotiny._0315_[30] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _09043_ (.RESET_B(net1570),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2025),
    .Q(\i_exotiny._0315_[31] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _09044_ (.RESET_B(net1359),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1206_ ),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r ),
    .CLK(clknet_5_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _09045_ (.RESET_B(net1358),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01102_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[0] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _09046_ (.RESET_B(net1356),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01103_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _09047_ (.RESET_B(net1571),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01104_),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _09048_ (.RESET_B(net804),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3391),
    .Q(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r [0]),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _09049_ (.RESET_B(net1354),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\i_exotiny._1266_ ),
    .Q(\i_exotiny._0352_ ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _09050_ (.RESET_B(net1352),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1884),
    .Q(\i_exotiny.i_rstctl.cnt[0] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _09051_ (.RESET_B(net1351),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01106_),
    .Q(\i_exotiny.i_rstctl.cnt[1] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _09052_ (.RESET_B(net1350),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2300),
    .Q(\i_exotiny.i_rstctl.cnt[2] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _09053_ (.RESET_B(net1349),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01108_),
    .Q(\i_exotiny.i_rstctl.cnt[3] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _09054_ (.RESET_B(net1348),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01109_),
    .Q(\i_exotiny.i_rstctl.cnt[4] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _09055_ (.RESET_B(net1347),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01110_),
    .Q(\i_exotiny.i_rstctl.cnt[5] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _09056_ (.RESET_B(net1346),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1971),
    .Q(\i_exotiny.i_rstctl.cnt[6] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _09057_ (.RESET_B(net1345),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01112_),
    .Q(\i_exotiny._1652_[0] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _09058_ (.RESET_B(net1344),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3725),
    .Q(\i_exotiny.i_wb_qspi_mem.cnt_r[1] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _09059_ (.RESET_B(net1343),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3701),
    .Q(\i_exotiny.i_wb_qspi_mem.cnt_r[2] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _09060_ (.RESET_B(net1342),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1831),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[0] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09061_ (.RESET_B(net1341),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01116_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[1] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09062_ (.RESET_B(net1340),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01117_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[2] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09063_ (.RESET_B(net1339),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1887),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[3] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09064_ (.RESET_B(net1338),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3629),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[4] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09065_ (.RESET_B(net1337),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01120_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[5] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _09066_ (.RESET_B(net1336),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1915),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[6] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _09067_ (.RESET_B(net1335),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2030),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[7] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _09068_ (.RESET_B(net1334),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01123_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[8] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _09069_ (.RESET_B(net1333),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01124_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[9] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09070_ (.RESET_B(net1332),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1879),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[10] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _09071_ (.RESET_B(net1331),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01126_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[11] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09072_ (.RESET_B(net1330),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1892),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[12] ),
    .CLK(clknet_5_11__leaf_clk_regs));
 sg13g2_dfrbpq_1 _09073_ (.RESET_B(net1329),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3237),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[13] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09074_ (.RESET_B(net1328),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01129_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[14] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09075_ (.RESET_B(net1327),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01130_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[15] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09076_ (.RESET_B(net1326),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1882),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[16] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09077_ (.RESET_B(net1325),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2056),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[17] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _09078_ (.RESET_B(net1324),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01133_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[18] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _09079_ (.RESET_B(net1323),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01134_),
    .Q(\i_exotiny.i_wdg_top.clk_div_inst.cnt[19] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_2 _09080_ (.RESET_B(net1322),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3106),
    .Q(\i_exotiny._0024_[0] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_2 _09081_ (.RESET_B(net1321),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2187),
    .Q(\i_exotiny._0024_[1] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_2 _09082_ (.RESET_B(net1320),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2463),
    .Q(\i_exotiny._0024_[2] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_2 _09083_ (.RESET_B(net1319),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2918),
    .Q(\i_exotiny._0024_[3] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09084_ (.RESET_B(net1318),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2098),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _09085_ (.RESET_B(net1317),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01140_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09086_ (.RESET_B(net1316),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01141_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _09087_ (.RESET_B(net1315),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2860),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _09088_ (.RESET_B(net1314),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01143_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _09089_ (.RESET_B(net1313),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01144_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09090_ (.RESET_B(net1312),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2687),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09091_ (.RESET_B(net1311),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2707),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _09092_ (.RESET_B(net1310),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01147_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _09093_ (.RESET_B(net1309),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01148_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09094_ (.RESET_B(net1308),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3339),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09095_ (.RESET_B(net1307),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01150_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09096_ (.RESET_B(net1306),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2786),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09097_ (.RESET_B(net1305),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3312),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09098_ (.RESET_B(net1304),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2131),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09099_ (.RESET_B(net1303),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01154_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _09100_ (.RESET_B(net1302),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2237),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09101_ (.RESET_B(net1301),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2397),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09102_ (.RESET_B(net1300),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01157_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09103_ (.RESET_B(net1299),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2350),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09104_ (.RESET_B(net1298),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01159_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _09105_ (.RESET_B(net1297),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01160_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09106_ (.RESET_B(net1296),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01161_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09107_ (.RESET_B(net1295),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01162_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _09108_ (.RESET_B(net1294),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3086),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _09109_ (.RESET_B(net1293),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01164_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _09110_ (.RESET_B(net1292),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2297),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _09111_ (.RESET_B(net871),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3146),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_2 _09112_ (.RESET_B(net870),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2183),
    .Q(\i_exotiny._0030_[0] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _09113_ (.RESET_B(net869),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01168_),
    .Q(\i_exotiny._0030_[1] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_2 _09114_ (.RESET_B(net868),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01169_),
    .Q(\i_exotiny._0030_[2] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _09115_ (.RESET_B(net867),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2634),
    .Q(\i_exotiny._0030_[3] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _09116_ (.RESET_B(net866),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01171_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09117_ (.RESET_B(net865),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01172_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09118_ (.RESET_B(net864),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01173_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _09119_ (.RESET_B(net863),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01174_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09120_ (.RESET_B(net862),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01175_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _09121_ (.RESET_B(net861),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2302),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09122_ (.RESET_B(net860),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01177_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09123_ (.RESET_B(net859),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01178_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09124_ (.RESET_B(net858),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2421),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _09125_ (.RESET_B(net857),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3139),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _09126_ (.RESET_B(net856),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3182),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _09127_ (.RESET_B(net855),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01182_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09128_ (.RESET_B(net854),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01183_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _09129_ (.RESET_B(net853),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2195),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _09130_ (.RESET_B(net852),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01185_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _09131_ (.RESET_B(net851),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2177),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _09132_ (.RESET_B(net850),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2527),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _09133_ (.RESET_B(net849),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01188_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _09134_ (.RESET_B(net848),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2500),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _09135_ (.RESET_B(net847),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01190_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _09136_ (.RESET_B(net846),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01191_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _09137_ (.RESET_B(net845),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2728),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _09138_ (.RESET_B(net844),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2173),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09139_ (.RESET_B(net843),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2210),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _09140_ (.RESET_B(net842),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2977),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _09141_ (.RESET_B(net841),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01196_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _09142_ (.RESET_B(net840),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01197_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _09143_ (.RESET_B(net839),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01198_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_2 _09144_ (.RESET_B(net838),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2993),
    .Q(\i_exotiny._0027_[0] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_2 _09145_ (.RESET_B(net837),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01200_),
    .Q(\i_exotiny._0027_[1] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_2 _09146_ (.RESET_B(net836),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01201_),
    .Q(\i_exotiny._0027_[2] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_2 _09147_ (.RESET_B(net835),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01202_),
    .Q(\i_exotiny._0027_[3] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _09148_ (.RESET_B(net834),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2991),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _09149_ (.RESET_B(net833),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01204_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _09150_ (.RESET_B(net832),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2725),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09151_ (.RESET_B(net831),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3177),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _09152_ (.RESET_B(net830),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2336),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _09153_ (.RESET_B(net829),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2546),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _09154_ (.RESET_B(net828),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3272),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09155_ (.RESET_B(net827),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01210_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _09156_ (.RESET_B(net826),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01211_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _09157_ (.RESET_B(net825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2580),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _09158_ (.RESET_B(net824),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2423),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09159_ (.RESET_B(net823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2569),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _09160_ (.RESET_B(net822),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01215_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _09161_ (.RESET_B(net821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01216_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _09162_ (.RESET_B(net820),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01217_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _09163_ (.RESET_B(net819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01218_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _09164_ (.RESET_B(net818),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2049),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _09165_ (.RESET_B(net817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2749),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _09166_ (.RESET_B(net816),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01221_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _09167_ (.RESET_B(net815),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2388),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _09168_ (.RESET_B(net814),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01223_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _09169_ (.RESET_B(net813),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2380),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _09170_ (.RESET_B(net812),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2518),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _09171_ (.RESET_B(net811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01226_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _09172_ (.RESET_B(net810),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01227_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _09173_ (.RESET_B(net809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01228_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _09174_ (.RESET_B(net808),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01229_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _09175_ (.RESET_B(net807),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01230_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _09176_ (.RESET_B(net806),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3806),
    .Q(\i_exotiny.i_wb_spi.sck_r ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _09177_ (.RESET_B(net805),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1962),
    .Q(\i_exotiny._1924_[1] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _09178_ (.RESET_B(net803),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3158),
    .Q(\i_exotiny._0026_[0] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _09179_ (.RESET_B(net802),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2601),
    .Q(\i_exotiny._0026_[1] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _09180_ (.RESET_B(net801),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01235_),
    .Q(\i_exotiny._0026_[2] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _09181_ (.RESET_B(net800),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01236_),
    .Q(\i_exotiny._0026_[3] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _09182_ (.RESET_B(net799),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01237_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09183_ (.RESET_B(net798),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01238_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _09184_ (.RESET_B(net797),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01239_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09185_ (.RESET_B(net796),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2461),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _09186_ (.RESET_B(net795),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2405),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09187_ (.RESET_B(net794),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2901),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _09188_ (.RESET_B(net793),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3058),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09189_ (.RESET_B(net792),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2744),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09190_ (.RESET_B(net791),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01245_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09191_ (.RESET_B(net790),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2242),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09192_ (.RESET_B(net789),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2582),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09193_ (.RESET_B(net788),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01248_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09194_ (.RESET_B(net787),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01249_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09195_ (.RESET_B(net786),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01250_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09196_ (.RESET_B(net785),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01251_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09197_ (.RESET_B(net784),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01252_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09198_ (.RESET_B(net783),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2838),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09199_ (.RESET_B(net782),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01254_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09200_ (.RESET_B(net781),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2133),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09201_ (.RESET_B(net780),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2520),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09202_ (.RESET_B(net779),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01257_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09203_ (.RESET_B(net778),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2697),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09204_ (.RESET_B(net777),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01259_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _09205_ (.RESET_B(net776),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2560),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _09206_ (.RESET_B(net773),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3008),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _09207_ (.RESET_B(net772),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3051),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _09208_ (.RESET_B(net771),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01263_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _09209_ (.RESET_B(net770),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2854),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _09210_ (.RESET_B(net769),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3228),
    .Q(\i_exotiny._0023_[0] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_2 _09211_ (.RESET_B(net768),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3204),
    .Q(\i_exotiny._0023_[1] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_2 _09212_ (.RESET_B(net767),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01267_),
    .Q(\i_exotiny._0023_[2] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_2 _09213_ (.RESET_B(net766),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01268_),
    .Q(\i_exotiny._0023_[3] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09214_ (.RESET_B(net765),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2072),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09215_ (.RESET_B(net764),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01270_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09216_ (.RESET_B(net763),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01271_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09217_ (.RESET_B(net762),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3293),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _09218_ (.RESET_B(net761),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01273_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09219_ (.RESET_B(net760),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2834),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09220_ (.RESET_B(net759),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01275_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09221_ (.RESET_B(net758),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2252),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _09222_ (.RESET_B(net757),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01277_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09223_ (.RESET_B(net756),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01278_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09224_ (.RESET_B(net755),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2752),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09225_ (.RESET_B(net754),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01280_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _09226_ (.RESET_B(net753),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2870),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09227_ (.RESET_B(net752),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2626),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09228_ (.RESET_B(net751),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01283_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09229_ (.RESET_B(net750),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2346),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _09230_ (.RESET_B(net749),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3226),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _09231_ (.RESET_B(net748),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01286_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09232_ (.RESET_B(net747),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01287_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09233_ (.RESET_B(net746),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01288_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _09234_ (.RESET_B(net745),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01289_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09235_ (.RESET_B(net744),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2681),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09236_ (.RESET_B(net704),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01291_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09237_ (.RESET_B(net701),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2498),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _09238_ (.RESET_B(net699),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3018),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09239_ (.RESET_B(net697),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3376),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09240_ (.RESET_B(net567),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2705),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _09241_ (.RESET_B(net566),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01296_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_2 _09242_ (.RESET_B(net565),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2135),
    .Q(\i_exotiny._0022_[0] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_2 _09243_ (.RESET_B(net564),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3492),
    .Q(\i_exotiny._0022_[1] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_2 _09244_ (.RESET_B(net563),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2163),
    .Q(\i_exotiny._0022_[2] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_2 _09245_ (.RESET_B(net562),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2308),
    .Q(\i_exotiny._0022_[3] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _09246_ (.RESET_B(net561),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01301_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09247_ (.RESET_B(net560),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3125),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09248_ (.RESET_B(net559),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01303_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _09249_ (.RESET_B(net558),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01304_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _09250_ (.RESET_B(net557),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01305_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09251_ (.RESET_B(net556),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01306_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09252_ (.RESET_B(net555),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2143),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09253_ (.RESET_B(net554),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01308_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09254_ (.RESET_B(net553),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2809),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09255_ (.RESET_B(net552),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01310_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09256_ (.RESET_B(net551),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01311_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09257_ (.RESET_B(net550),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01312_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09258_ (.RESET_B(net509),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01313_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09259_ (.RESET_B(net243),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01314_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09260_ (.RESET_B(net241),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2923),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _09261_ (.RESET_B(net239),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3421),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _09262_ (.RESET_B(net237),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2470),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09263_ (.RESET_B(net235),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2348),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _09264_ (.RESET_B(net101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3253),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09265_ (.RESET_B(net99),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2537),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09266_ (.RESET_B(net97),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01321_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09267_ (.RESET_B(net93),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01322_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09268_ (.RESET_B(net91),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2122),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09269_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2268),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _09270_ (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2472),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09271_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2911),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _09272_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01327_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _09273_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01328_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _09274_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2070),
    .Q(\i_exotiny._0021_[0] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_2 _09275_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2372),
    .Q(\i_exotiny._0021_[1] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_2 _09276_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2452),
    .Q(\i_exotiny._0021_[2] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_2 _09277_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01332_),
    .Q(\i_exotiny._0021_[3] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _09278_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01333_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[4] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _09279_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2366),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[5] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _09280_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01335_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[6] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _09281_ (.RESET_B(net59),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3141),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[7] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _09282_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2685),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[8] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _09283_ (.RESET_B(net55),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01338_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[9] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _09284_ (.RESET_B(net53),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01339_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[10] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _09285_ (.RESET_B(net51),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2189),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[11] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _09286_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3474),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[12] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _09287_ (.RESET_B(net1825),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2212),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[13] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _09288_ (.RESET_B(net1823),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3251),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[14] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _09289_ (.RESET_B(net1821),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01344_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[15] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _09290_ (.RESET_B(net1819),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2328),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[16] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _09291_ (.RESET_B(net1817),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01346_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[17] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _09292_ (.RESET_B(net1815),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2260),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[18] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _09293_ (.RESET_B(net1813),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01348_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[19] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09294_ (.RESET_B(net1811),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01349_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[20] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _09295_ (.RESET_B(net1809),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01350_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[21] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _09296_ (.RESET_B(net1771),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01351_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[22] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _09297_ (.RESET_B(net1769),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2191),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[23] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _09298_ (.RESET_B(net1767),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2254),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[24] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _09299_ (.RESET_B(net1539),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net2811),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[25] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _09300_ (.RESET_B(net1537),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01355_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[26] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _09301_ (.RESET_B(net1535),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01356_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[27] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _09302_ (.RESET_B(net1533),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01357_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[28] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _09303_ (.RESET_B(net1357),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3098),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[29] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _09304_ (.RESET_B(net1355),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net3067),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[30] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _09305_ (.RESET_B(net1353),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01360_),
    .Q(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[31] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_tiehi _07904__43 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net43));
 sg13g2_tiehi _07898__44 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net44));
 sg13g2_tiehi _07899__45 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net45));
 sg13g2_tiehi _07900__46 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net46));
 sg13g2_tiehi _07901__47 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net47));
 sg13g2_tiehi _07902__48 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net48));
 sg13g2_tiehi _08577__49 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net49));
 sg13g2_tiehi _07903__50 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net50));
 sg13g2_tiehi _09285__51 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net51));
 sg13g2_tiehi _08576__52 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net52));
 sg13g2_tiehi _09284__53 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net53));
 sg13g2_tiehi _08575__54 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net54));
 sg13g2_tiehi _09283__55 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net55));
 sg13g2_tiehi _08574__56 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net56));
 sg13g2_tiehi _09282__57 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net57));
 sg13g2_tiehi _08573__58 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net58));
 sg13g2_tiehi _09281__59 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net59));
 sg13g2_tiehi _08572__60 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net60));
 sg13g2_tiehi _09280__61 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net61));
 sg13g2_tiehi _08571__62 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net62));
 sg13g2_tiehi _09279__63 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net63));
 sg13g2_tiehi _08570__64 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net64));
 sg13g2_tiehi _09278__65 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net65));
 sg13g2_tiehi _08569__66 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net66));
 sg13g2_tiehi _09277__67 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net67));
 sg13g2_tiehi _08568__68 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net68));
 sg13g2_tiehi _09276__69 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net69));
 sg13g2_tiehi _08567__70 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net70));
 sg13g2_tiehi _09275__71 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net71));
 sg13g2_tiehi _08566__72 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net72));
 sg13g2_tiehi _09274__73 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net73));
 sg13g2_tiehi _08565__74 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net74));
 sg13g2_tiehi _09273__75 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net75));
 sg13g2_tiehi _08564__76 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net76));
 sg13g2_tiehi _09272__77 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net77));
 sg13g2_tiehi _08563__78 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net78));
 sg13g2_tiehi _09271__79 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net79));
 sg13g2_tiehi _08562__80 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net80));
 sg13g2_tiehi _09270__81 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net81));
 sg13g2_tiehi _08561__82 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net82));
 sg13g2_tiehi _09269__83 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net83));
 sg13g2_tiehi _08560__84 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net84));
 sg13g2_tiehi _07941__85 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net85));
 sg13g2_tiehi _07942__86 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net86));
 sg13g2_tiehi _07943__87 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net87));
 sg13g2_tiehi _07944__88 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net88));
 sg13g2_tiehi _07945__89 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net89));
 sg13g2_tiehi _07946__90 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net90));
 sg13g2_tiehi _09268__91 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net91));
 sg13g2_tiehi _08559__92 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net92));
 sg13g2_tiehi _09267__93 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net93));
 sg13g2_tiehi _07947__94 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net94));
 sg13g2_tiehi _07951__95 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net95));
 sg13g2_tiehi _08558__96 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net96));
 sg13g2_tiehi _09266__97 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net97));
 sg13g2_tiehi _08557__98 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net98));
 sg13g2_tiehi _09265__99 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net99));
 sg13g2_tiehi _08556__100 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net100));
 sg13g2_tiehi _09264__101 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net101));
 sg13g2_tiehi _08555__102 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net102));
 sg13g2_tiehi _08554__103 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net103));
 sg13g2_tiehi _08552__104 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net104));
 sg13g2_tiehi _08551__105 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net105));
 sg13g2_tiehi _08550__106 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net106));
 sg13g2_tiehi _08549__107 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net107));
 sg13g2_tiehi _08548__108 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net108));
 sg13g2_tiehi _08547__109 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net109));
 sg13g2_tiehi _08546__110 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net110));
 sg13g2_tiehi _08545__111 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net111));
 sg13g2_tiehi _08544__112 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net112));
 sg13g2_tiehi _08543__113 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net113));
 sg13g2_tiehi _07973__114 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net114));
 sg13g2_tiehi _07974__115 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net115));
 sg13g2_tiehi _07975__116 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net116));
 sg13g2_tiehi _07976__117 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net117));
 sg13g2_tiehi _07977__118 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net118));
 sg13g2_tiehi _07978__119 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net119));
 sg13g2_tiehi _07979__120 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net120));
 sg13g2_tiehi _07980__121 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net121));
 sg13g2_tiehi _07981__122 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net122));
 sg13g2_tiehi _07982__123 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net123));
 sg13g2_tiehi _07983__124 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net124));
 sg13g2_tiehi _07984__125 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net125));
 sg13g2_tiehi _07985__126 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net126));
 sg13g2_tiehi _07986__127 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net127));
 sg13g2_tiehi _07987__128 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net128));
 sg13g2_tiehi _07988__129 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net129));
 sg13g2_tiehi _07989__130 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net130));
 sg13g2_tiehi _07990__131 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net131));
 sg13g2_tiehi _07991__132 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net132));
 sg13g2_tiehi _07992__133 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net133));
 sg13g2_tiehi _07993__134 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net134));
 sg13g2_tiehi _07994__135 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net135));
 sg13g2_tiehi _07995__136 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net136));
 sg13g2_tiehi _07996__137 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net137));
 sg13g2_tiehi _08542__138 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net138));
 sg13g2_tiehi _08541__139 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net139));
 sg13g2_tiehi _08540__140 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net140));
 sg13g2_tiehi _08539__141 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net141));
 sg13g2_tiehi _08538__142 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net142));
 sg13g2_tiehi _08537__143 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net143));
 sg13g2_tiehi _08536__144 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net144));
 sg13g2_tiehi _08535__145 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net145));
 sg13g2_tiehi _08534__146 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net146));
 sg13g2_tiehi _08533__147 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net147));
 sg13g2_tiehi _08532__148 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net148));
 sg13g2_tiehi _08531__149 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net149));
 sg13g2_tiehi _08530__150 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net150));
 sg13g2_tiehi _08529__151 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net151));
 sg13g2_tiehi _08528__152 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net152));
 sg13g2_tiehi _08527__153 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net153));
 sg13g2_tiehi _08526__154 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net154));
 sg13g2_tiehi _08525__155 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net155));
 sg13g2_tiehi _08524__156 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net156));
 sg13g2_tiehi _08523__157 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net157));
 sg13g2_tiehi _08522__158 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net158));
 sg13g2_tiehi _08521__159 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net159));
 sg13g2_tiehi _08520__160 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net160));
 sg13g2_tiehi _08519__161 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net161));
 sg13g2_tiehi _08518__162 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net162));
 sg13g2_tiehi _08517__163 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net163));
 sg13g2_tiehi _08516__164 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net164));
 sg13g2_tiehi _08515__165 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net165));
 sg13g2_tiehi _08514__166 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net166));
 sg13g2_tiehi _08513__167 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net167));
 sg13g2_tiehi _08512__168 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net168));
 sg13g2_tiehi _08511__169 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net169));
 sg13g2_tiehi _08510__170 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net170));
 sg13g2_tiehi _08509__171 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net171));
 sg13g2_tiehi _08508__172 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net172));
 sg13g2_tiehi _08507__173 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net173));
 sg13g2_tiehi _08506__174 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net174));
 sg13g2_tiehi _08505__175 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net175));
 sg13g2_tiehi _08504__176 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net176));
 sg13g2_tiehi _08503__177 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net177));
 sg13g2_tiehi _08502__178 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net178));
 sg13g2_tiehi _08501__179 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net179));
 sg13g2_tiehi _08500__180 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net180));
 sg13g2_tiehi _08499__181 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net181));
 sg13g2_tiehi _08498__182 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net182));
 sg13g2_tiehi _08497__183 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net183));
 sg13g2_tiehi _08496__184 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net184));
 sg13g2_tiehi _08495__185 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net185));
 sg13g2_tiehi _08494__186 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net186));
 sg13g2_tiehi _08493__187 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net187));
 sg13g2_tiehi _08492__188 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net188));
 sg13g2_tiehi _08491__189 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net189));
 sg13g2_tiehi _08490__190 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net190));
 sg13g2_tiehi _08489__191 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net191));
 sg13g2_tiehi _08488__192 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net192));
 sg13g2_tiehi _08487__193 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net193));
 sg13g2_tiehi _08486__194 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net194));
 sg13g2_tiehi _08485__195 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net195));
 sg13g2_tiehi _08484__196 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net196));
 sg13g2_tiehi _08483__197 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net197));
 sg13g2_tiehi _08482__198 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net198));
 sg13g2_tiehi _08481__199 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net199));
 sg13g2_tiehi _08480__200 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net200));
 sg13g2_tiehi _08479__201 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net201));
 sg13g2_tiehi _08478__202 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net202));
 sg13g2_tiehi _08477__203 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net203));
 sg13g2_tiehi _08476__204 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net204));
 sg13g2_tiehi _08475__205 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net205));
 sg13g2_tiehi _08474__206 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net206));
 sg13g2_tiehi _08473__207 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net207));
 sg13g2_tiehi _08472__208 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net208));
 sg13g2_tiehi _08471__209 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net209));
 sg13g2_tiehi _08470__210 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net210));
 sg13g2_tiehi _08469__211 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net211));
 sg13g2_tiehi _08468__212 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net212));
 sg13g2_tiehi _08467__213 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net213));
 sg13g2_tiehi _08466__214 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net214));
 sg13g2_tiehi _08465__215 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net215));
 sg13g2_tiehi _08464__216 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net216));
 sg13g2_tiehi _08463__217 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net217));
 sg13g2_tiehi _08462__218 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net218));
 sg13g2_tiehi _08461__219 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net219));
 sg13g2_tiehi _08460__220 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net220));
 sg13g2_tiehi _08459__221 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net221));
 sg13g2_tiehi _08458__222 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net222));
 sg13g2_tiehi _08457__223 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net223));
 sg13g2_tiehi _08456__224 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net224));
 sg13g2_tiehi _08455__225 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net225));
 sg13g2_tiehi _08454__226 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net226));
 sg13g2_tiehi _08453__227 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net227));
 sg13g2_tiehi _08452__228 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net228));
 sg13g2_tiehi _08451__229 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net229));
 sg13g2_tiehi _08450__230 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net230));
 sg13g2_tiehi _08449__231 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net231));
 sg13g2_tiehi _08448__232 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net232));
 sg13g2_tiehi _08447__233 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net233));
 sg13g2_tiehi _08446__234 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net234));
 sg13g2_tiehi _09263__235 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net235));
 sg13g2_tiehi _08445__236 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net236));
 sg13g2_tiehi _09262__237 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net237));
 sg13g2_tiehi _08444__238 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net238));
 sg13g2_tiehi _09261__239 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net239));
 sg13g2_tiehi _08443__240 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net240));
 sg13g2_tiehi _09260__241 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net241));
 sg13g2_tiehi _08442__242 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net242));
 sg13g2_tiehi _09259__243 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net243));
 sg13g2_tiehi _08441__244 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net244));
 sg13g2_tiehi _08440__245 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net245));
 sg13g2_tiehi _08439__246 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net246));
 sg13g2_tiehi _08438__247 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net247));
 sg13g2_tiehi _08437__248 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net248));
 sg13g2_tiehi _08436__249 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net249));
 sg13g2_tiehi _08435__250 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net250));
 sg13g2_tiehi _08434__251 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net251));
 sg13g2_tiehi _08433__252 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net252));
 sg13g2_tiehi _08432__253 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net253));
 sg13g2_tiehi _08431__254 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net254));
 sg13g2_tiehi _08430__255 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net255));
 sg13g2_tiehi _08429__256 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net256));
 sg13g2_tiehi _08428__257 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net257));
 sg13g2_tiehi _08427__258 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net258));
 sg13g2_tiehi _08426__259 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net259));
 sg13g2_tiehi _08425__260 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net260));
 sg13g2_tiehi _08424__261 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net261));
 sg13g2_tiehi _08423__262 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net262));
 sg13g2_tiehi _08422__263 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net263));
 sg13g2_tiehi _08421__264 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net264));
 sg13g2_tiehi _08420__265 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net265));
 sg13g2_tiehi _08419__266 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net266));
 sg13g2_tiehi _08418__267 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net267));
 sg13g2_tiehi _08417__268 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net268));
 sg13g2_tiehi _08416__269 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net269));
 sg13g2_tiehi _08415__270 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net270));
 sg13g2_tiehi _08414__271 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net271));
 sg13g2_tiehi _08413__272 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net272));
 sg13g2_tiehi _08412__273 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net273));
 sg13g2_tiehi _08411__274 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net274));
 sg13g2_tiehi _08410__275 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net275));
 sg13g2_tiehi _08409__276 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net276));
 sg13g2_tiehi _08408__277 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net277));
 sg13g2_tiehi _08407__278 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net278));
 sg13g2_tiehi _08406__279 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net279));
 sg13g2_tiehi _08405__280 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net280));
 sg13g2_tiehi _08404__281 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net281));
 sg13g2_tiehi _08403__282 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net282));
 sg13g2_tiehi _08402__283 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net283));
 sg13g2_tiehi _08401__284 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net284));
 sg13g2_tiehi _08400__285 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net285));
 sg13g2_tiehi _08392__286 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net286));
 sg13g2_tiehi _08391__287 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net287));
 sg13g2_tiehi _08390__288 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net288));
 sg13g2_tiehi _08389__289 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net289));
 sg13g2_tiehi _08388__290 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net290));
 sg13g2_tiehi _08387__291 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net291));
 sg13g2_tiehi _08386__292 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net292));
 sg13g2_tiehi _08385__293 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net293));
 sg13g2_tiehi _08384__294 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net294));
 sg13g2_tiehi _08383__295 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net295));
 sg13g2_tiehi _08382__296 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net296));
 sg13g2_tiehi _08381__297 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net297));
 sg13g2_tiehi _08380__298 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net298));
 sg13g2_tiehi _08379__299 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net299));
 sg13g2_tiehi _08378__300 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net300));
 sg13g2_tiehi _08377__301 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net301));
 sg13g2_tiehi _08376__302 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net302));
 sg13g2_tiehi _08375__303 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net303));
 sg13g2_tiehi _08374__304 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net304));
 sg13g2_tiehi _08373__305 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net305));
 sg13g2_tiehi _08372__306 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net306));
 sg13g2_tiehi _08371__307 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net307));
 sg13g2_tiehi _08370__308 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net308));
 sg13g2_tiehi _08369__309 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net309));
 sg13g2_tiehi _08368__310 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net310));
 sg13g2_tiehi _08367__311 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net311));
 sg13g2_tiehi _08366__312 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net312));
 sg13g2_tiehi _08365__313 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net313));
 sg13g2_tiehi _08364__314 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net314));
 sg13g2_tiehi _08363__315 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net315));
 sg13g2_tiehi _08362__316 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net316));
 sg13g2_tiehi _08361__317 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net317));
 sg13g2_tiehi _08360__318 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net318));
 sg13g2_tiehi _08359__319 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net319));
 sg13g2_tiehi _08358__320 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net320));
 sg13g2_tiehi _08357__321 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net321));
 sg13g2_tiehi _08356__322 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net322));
 sg13g2_tiehi _08355__323 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net323));
 sg13g2_tiehi _08354__324 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net324));
 sg13g2_tiehi _08353__325 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net325));
 sg13g2_tiehi _08352__326 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net326));
 sg13g2_tiehi _08351__327 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net327));
 sg13g2_tiehi _08350__328 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net328));
 sg13g2_tiehi _08349__329 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net329));
 sg13g2_tiehi _08348__330 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net330));
 sg13g2_tiehi _08347__331 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net331));
 sg13g2_tiehi _08346__332 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net332));
 sg13g2_tiehi _08345__333 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net333));
 sg13g2_tiehi _08344__334 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net334));
 sg13g2_tiehi _08343__335 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net335));
 sg13g2_tiehi _08342__336 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net336));
 sg13g2_tiehi _08341__337 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net337));
 sg13g2_tiehi _08340__338 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net338));
 sg13g2_tiehi _08339__339 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net339));
 sg13g2_tiehi _08338__340 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net340));
 sg13g2_tiehi _08337__341 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net341));
 sg13g2_tiehi _08336__342 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net342));
 sg13g2_tiehi _08335__343 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net343));
 sg13g2_tiehi _08334__344 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net344));
 sg13g2_tiehi _08333__345 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net345));
 sg13g2_tiehi _08332__346 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net346));
 sg13g2_tiehi _08331__347 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net347));
 sg13g2_tiehi _08330__348 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net348));
 sg13g2_tiehi _08329__349 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net349));
 sg13g2_tiehi _08328__350 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net350));
 sg13g2_tiehi _08327__351 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net351));
 sg13g2_tiehi _08326__352 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net352));
 sg13g2_tiehi _08325__353 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net353));
 sg13g2_tiehi _08324__354 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net354));
 sg13g2_tiehi _08323__355 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net355));
 sg13g2_tiehi _08322__356 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net356));
 sg13g2_tiehi _08321__357 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net357));
 sg13g2_tiehi _08320__358 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net358));
 sg13g2_tiehi _08319__359 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net359));
 sg13g2_tiehi _08318__360 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net360));
 sg13g2_tiehi _08317__361 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net361));
 sg13g2_tiehi _08316__362 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net362));
 sg13g2_tiehi _08315__363 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net363));
 sg13g2_tiehi _08314__364 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net364));
 sg13g2_tiehi _08313__365 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net365));
 sg13g2_tiehi _08312__366 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net366));
 sg13g2_tiehi _08311__367 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net367));
 sg13g2_tiehi _08310__368 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net368));
 sg13g2_tiehi _08309__369 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net369));
 sg13g2_tiehi _08308__370 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net370));
 sg13g2_tiehi _08307__371 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net371));
 sg13g2_tiehi _08306__372 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net372));
 sg13g2_tiehi _08305__373 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net373));
 sg13g2_tiehi _08304__374 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net374));
 sg13g2_tiehi _08303__375 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net375));
 sg13g2_tiehi _08302__376 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net376));
 sg13g2_tiehi _08301__377 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net377));
 sg13g2_tiehi _08300__378 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net378));
 sg13g2_tiehi _08299__379 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net379));
 sg13g2_tiehi _08298__380 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net380));
 sg13g2_tiehi _08297__381 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net381));
 sg13g2_tiehi _08296__382 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net382));
 sg13g2_tiehi _08295__383 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net383));
 sg13g2_tiehi _08294__384 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net384));
 sg13g2_tiehi _08293__385 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net385));
 sg13g2_tiehi _08292__386 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net386));
 sg13g2_tiehi _08291__387 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net387));
 sg13g2_tiehi _08290__388 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net388));
 sg13g2_tiehi _08289__389 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net389));
 sg13g2_tiehi _08288__390 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net390));
 sg13g2_tiehi _08287__391 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net391));
 sg13g2_tiehi _08286__392 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net392));
 sg13g2_tiehi _08285__393 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net393));
 sg13g2_tiehi _08284__394 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net394));
 sg13g2_tiehi _08283__395 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net395));
 sg13g2_tiehi _08282__396 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net396));
 sg13g2_tiehi _08281__397 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net397));
 sg13g2_tiehi _08280__398 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net398));
 sg13g2_tiehi _08279__399 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net399));
 sg13g2_tiehi _08278__400 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net400));
 sg13g2_tiehi _08277__401 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net401));
 sg13g2_tiehi _08276__402 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net402));
 sg13g2_tiehi _08275__403 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net403));
 sg13g2_tiehi _08274__404 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net404));
 sg13g2_tiehi _08273__405 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net405));
 sg13g2_tiehi _08272__406 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net406));
 sg13g2_tiehi _08271__407 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net407));
 sg13g2_tiehi _08270__408 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net408));
 sg13g2_tiehi _08269__409 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net409));
 sg13g2_tiehi _08268__410 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net410));
 sg13g2_tiehi _08267__411 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net411));
 sg13g2_tiehi _08266__412 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net412));
 sg13g2_tiehi _08264__413 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net413));
 sg13g2_tiehi _08263__414 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net414));
 sg13g2_tiehi _08262__415 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net415));
 sg13g2_tiehi _08261__416 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net416));
 sg13g2_tiehi _08260__417 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net417));
 sg13g2_tiehi _08259__418 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net418));
 sg13g2_tiehi _08258__419 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net419));
 sg13g2_tiehi _08257__420 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net420));
 sg13g2_tiehi _08256__421 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net421));
 sg13g2_tiehi _08255__422 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net422));
 sg13g2_tiehi _08254__423 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net423));
 sg13g2_tiehi _08253__424 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net424));
 sg13g2_tiehi _08252__425 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net425));
 sg13g2_tiehi _08251__426 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net426));
 sg13g2_tiehi _08250__427 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net427));
 sg13g2_tiehi _08249__428 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net428));
 sg13g2_tiehi _08248__429 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net429));
 sg13g2_tiehi _08247__430 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net430));
 sg13g2_tiehi _08246__431 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net431));
 sg13g2_tiehi _08245__432 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net432));
 sg13g2_tiehi _08244__433 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net433));
 sg13g2_tiehi _08243__434 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net434));
 sg13g2_tiehi _08242__435 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net435));
 sg13g2_tiehi _08241__436 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net436));
 sg13g2_tiehi _08240__437 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net437));
 sg13g2_tiehi _08239__438 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net438));
 sg13g2_tiehi _08238__439 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net439));
 sg13g2_tiehi _08237__440 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net440));
 sg13g2_tiehi _08236__441 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net441));
 sg13g2_tiehi _08235__442 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net442));
 sg13g2_tiehi _08234__443 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net443));
 sg13g2_tiehi _08233__444 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net444));
 sg13g2_tiehi _08232__445 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net445));
 sg13g2_tiehi _08231__446 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net446));
 sg13g2_tiehi _08230__447 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net447));
 sg13g2_tiehi _08229__448 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net448));
 sg13g2_tiehi _08228__449 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net449));
 sg13g2_tiehi _08227__450 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net450));
 sg13g2_tiehi _08226__451 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net451));
 sg13g2_tiehi _08225__452 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net452));
 sg13g2_tiehi _08224__453 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net453));
 sg13g2_tiehi _08223__454 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net454));
 sg13g2_tiehi _08222__455 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net455));
 sg13g2_tiehi _08221__456 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net456));
 sg13g2_tiehi _08220__457 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net457));
 sg13g2_tiehi _08219__458 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net458));
 sg13g2_tiehi _08218__459 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net459));
 sg13g2_tiehi _08217__460 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net460));
 sg13g2_tiehi _08216__461 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net461));
 sg13g2_tiehi _08215__462 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net462));
 sg13g2_tiehi _08214__463 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net463));
 sg13g2_tiehi _08213__464 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net464));
 sg13g2_tiehi _08212__465 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net465));
 sg13g2_tiehi _08211__466 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net466));
 sg13g2_tiehi _08210__467 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net467));
 sg13g2_tiehi _08209__468 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net468));
 sg13g2_tiehi _08208__469 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net469));
 sg13g2_tiehi _08207__470 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net470));
 sg13g2_tiehi _08206__471 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net471));
 sg13g2_tiehi _08205__472 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net472));
 sg13g2_tiehi _08204__473 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net473));
 sg13g2_tiehi _08203__474 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net474));
 sg13g2_tiehi _08202__475 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net475));
 sg13g2_tiehi _08201__476 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net476));
 sg13g2_tiehi _08200__477 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net477));
 sg13g2_tiehi _08199__478 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net478));
 sg13g2_tiehi _08198__479 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net479));
 sg13g2_tiehi _08197__480 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net480));
 sg13g2_tiehi _08196__481 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net481));
 sg13g2_tiehi _08195__482 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net482));
 sg13g2_tiehi _08194__483 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net483));
 sg13g2_tiehi _08193__484 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net484));
 sg13g2_tiehi _08192__485 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net485));
 sg13g2_tiehi _08191__486 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net486));
 sg13g2_tiehi _08190__487 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net487));
 sg13g2_tiehi _08189__488 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net488));
 sg13g2_tiehi _08188__489 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net489));
 sg13g2_tiehi _08187__490 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net490));
 sg13g2_tiehi _08186__491 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net491));
 sg13g2_tiehi _08185__492 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net492));
 sg13g2_tiehi _08184__493 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net493));
 sg13g2_tiehi _08183__494 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net494));
 sg13g2_tiehi _08182__495 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net495));
 sg13g2_tiehi _08181__496 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net496));
 sg13g2_tiehi _08180__497 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net497));
 sg13g2_tiehi _08179__498 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net498));
 sg13g2_tiehi _08178__499 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net499));
 sg13g2_tiehi _08177__500 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net500));
 sg13g2_tiehi _08176__501 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net501));
 sg13g2_tiehi _08175__502 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net502));
 sg13g2_tiehi _08174__503 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net503));
 sg13g2_tiehi _08173__504 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net504));
 sg13g2_tiehi _08172__505 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net505));
 sg13g2_tiehi _08171__506 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net506));
 sg13g2_tiehi _08170__507 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net507));
 sg13g2_tiehi _08169__508 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net508));
 sg13g2_tiehi _09258__509 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net509));
 sg13g2_tiehi _08168__510 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net510));
 sg13g2_tiehi _08167__511 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net511));
 sg13g2_tiehi _08166__512 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net512));
 sg13g2_tiehi _08165__513 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net513));
 sg13g2_tiehi _08164__514 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net514));
 sg13g2_tiehi _08163__515 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net515));
 sg13g2_tiehi _08162__516 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net516));
 sg13g2_tiehi _08161__517 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net517));
 sg13g2_tiehi _08160__518 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net518));
 sg13g2_tiehi _08159__519 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net519));
 sg13g2_tiehi _08158__520 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net520));
 sg13g2_tiehi _08157__521 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net521));
 sg13g2_tiehi _08156__522 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net522));
 sg13g2_tiehi _08155__523 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net523));
 sg13g2_tiehi _08154__524 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net524));
 sg13g2_tiehi _08153__525 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net525));
 sg13g2_tiehi _08152__526 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net526));
 sg13g2_tiehi _08151__527 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net527));
 sg13g2_tiehi _08150__528 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net528));
 sg13g2_tiehi _08149__529 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net529));
 sg13g2_tiehi _08148__530 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net530));
 sg13g2_tiehi _08147__531 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net531));
 sg13g2_tiehi _07997__532 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net532));
 sg13g2_tiehi _08393__533 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net533));
 sg13g2_tiehi _08394__534 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net534));
 sg13g2_tiehi _08395__535 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net535));
 sg13g2_tiehi _08396__536 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net536));
 sg13g2_tiehi _08397__537 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net537));
 sg13g2_tiehi _08398__538 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net538));
 sg13g2_tiehi _08146__539 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net539));
 sg13g2_tiehi _08145__540 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net540));
 sg13g2_tiehi _08144__541 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net541));
 sg13g2_tiehi _08143__542 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net542));
 sg13g2_tiehi _08142__543 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net543));
 sg13g2_tiehi _08141__544 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net544));
 sg13g2_tiehi _08140__545 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net545));
 sg13g2_tiehi _08139__546 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net546));
 sg13g2_tiehi _08138__547 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net547));
 sg13g2_tiehi _08137__548 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net548));
 sg13g2_tiehi _08136__549 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net549));
 sg13g2_tiehi _09257__550 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net550));
 sg13g2_tiehi _09256__551 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net551));
 sg13g2_tiehi _09255__552 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net552));
 sg13g2_tiehi _09254__553 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net553));
 sg13g2_tiehi _09253__554 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net554));
 sg13g2_tiehi _09252__555 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net555));
 sg13g2_tiehi _09251__556 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net556));
 sg13g2_tiehi _09250__557 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net557));
 sg13g2_tiehi _09249__558 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net558));
 sg13g2_tiehi _09248__559 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net559));
 sg13g2_tiehi _09247__560 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net560));
 sg13g2_tiehi _09246__561 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net561));
 sg13g2_tiehi _09245__562 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net562));
 sg13g2_tiehi _09244__563 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net563));
 sg13g2_tiehi _09243__564 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net564));
 sg13g2_tiehi _09242__565 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net565));
 sg13g2_tiehi _09241__566 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net566));
 sg13g2_tiehi _09240__567 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net567));
 sg13g2_tiehi _08126__568 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net568));
 sg13g2_tiehi _08125__569 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net569));
 sg13g2_tiehi _08124__570 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net570));
 sg13g2_tiehi _08123__571 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net571));
 sg13g2_tiehi _08122__572 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net572));
 sg13g2_tiehi _08121__573 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net573));
 sg13g2_tiehi _08120__574 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net574));
 sg13g2_tiehi _08119__575 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net575));
 sg13g2_tiehi _08118__576 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net576));
 sg13g2_tiehi _08117__577 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net577));
 sg13g2_tiehi _08116__578 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net578));
 sg13g2_tiehi _08115__579 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net579));
 sg13g2_tiehi _08114__580 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net580));
 sg13g2_tiehi _08113__581 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net581));
 sg13g2_tiehi _08112__582 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net582));
 sg13g2_tiehi _08111__583 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net583));
 sg13g2_tiehi _08110__584 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net584));
 sg13g2_tiehi _08109__585 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net585));
 sg13g2_tiehi _08108__586 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net586));
 sg13g2_tiehi _08107__587 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net587));
 sg13g2_tiehi _08106__588 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net588));
 sg13g2_tiehi _08105__589 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net589));
 sg13g2_tiehi _08104__590 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net590));
 sg13g2_tiehi _08103__591 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net591));
 sg13g2_tiehi _08102__592 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net592));
 sg13g2_tiehi _08101__593 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net593));
 sg13g2_tiehi _08100__594 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net594));
 sg13g2_tiehi _08099__595 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net595));
 sg13g2_tiehi _08098__596 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net596));
 sg13g2_tiehi _08097__597 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net597));
 sg13g2_tiehi _08096__598 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net598));
 sg13g2_tiehi _08095__599 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net599));
 sg13g2_tiehi _08094__600 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net600));
 sg13g2_tiehi _08093__601 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net601));
 sg13g2_tiehi _08092__602 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net602));
 sg13g2_tiehi _08091__603 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net603));
 sg13g2_tiehi _08090__604 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net604));
 sg13g2_tiehi _08089__605 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net605));
 sg13g2_tiehi _08088__606 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net606));
 sg13g2_tiehi _08087__607 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net607));
 sg13g2_tiehi _08086__608 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net608));
 sg13g2_tiehi _08085__609 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net609));
 sg13g2_tiehi _08084__610 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net610));
 sg13g2_tiehi _08083__611 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net611));
 sg13g2_tiehi _08082__612 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net612));
 sg13g2_tiehi _08081__613 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net613));
 sg13g2_tiehi _08080__614 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net614));
 sg13g2_tiehi _08079__615 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net615));
 sg13g2_tiehi _08078__616 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net616));
 sg13g2_tiehi _08077__617 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net617));
 sg13g2_tiehi _08076__618 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net618));
 sg13g2_tiehi _08075__619 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net619));
 sg13g2_tiehi _08074__620 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net620));
 sg13g2_tiehi _08073__621 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net621));
 sg13g2_tiehi _08072__622 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net622));
 sg13g2_tiehi _08071__623 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net623));
 sg13g2_tiehi _08070__624 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net624));
 sg13g2_tiehi _08069__625 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net625));
 sg13g2_tiehi _08068__626 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net626));
 sg13g2_tiehi _08067__627 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net627));
 sg13g2_tiehi _08066__628 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net628));
 sg13g2_tiehi _08065__629 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net629));
 sg13g2_tiehi _08064__630 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net630));
 sg13g2_tiehi _08063__631 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net631));
 sg13g2_tiehi _08062__632 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net632));
 sg13g2_tiehi _08061__633 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net633));
 sg13g2_tiehi _08060__634 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net634));
 sg13g2_tiehi _08059__635 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net635));
 sg13g2_tiehi _08058__636 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net636));
 sg13g2_tiehi _08057__637 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net637));
 sg13g2_tiehi _08056__638 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net638));
 sg13g2_tiehi _08055__639 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net639));
 sg13g2_tiehi _08054__640 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net640));
 sg13g2_tiehi _08053__641 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net641));
 sg13g2_tiehi _08052__642 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net642));
 sg13g2_tiehi _08051__643 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net643));
 sg13g2_tiehi _08050__644 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net644));
 sg13g2_tiehi _08049__645 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net645));
 sg13g2_tiehi _08048__646 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net646));
 sg13g2_tiehi _08047__647 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net647));
 sg13g2_tiehi _08046__648 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net648));
 sg13g2_tiehi _08045__649 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net649));
 sg13g2_tiehi _08044__650 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net650));
 sg13g2_tiehi _08043__651 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net651));
 sg13g2_tiehi _08042__652 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net652));
 sg13g2_tiehi _08041__653 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net653));
 sg13g2_tiehi _08040__654 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net654));
 sg13g2_tiehi _08039__655 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net655));
 sg13g2_tiehi _08038__656 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net656));
 sg13g2_tiehi _08037__657 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net657));
 sg13g2_tiehi _08036__658 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net658));
 sg13g2_tiehi _08035__659 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net659));
 sg13g2_tiehi _08034__660 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net660));
 sg13g2_tiehi _08033__661 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net661));
 sg13g2_tiehi _08032__662 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net662));
 sg13g2_tiehi _08031__663 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net663));
 sg13g2_tiehi _08030__664 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net664));
 sg13g2_tiehi _08029__665 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net665));
 sg13g2_tiehi _08028__666 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net666));
 sg13g2_tiehi _08027__667 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net667));
 sg13g2_tiehi _08026__668 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net668));
 sg13g2_tiehi _08025__669 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net669));
 sg13g2_tiehi _08024__670 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net670));
 sg13g2_tiehi _08023__671 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net671));
 sg13g2_tiehi _08022__672 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net672));
 sg13g2_tiehi _08021__673 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net673));
 sg13g2_tiehi _08020__674 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net674));
 sg13g2_tiehi _08019__675 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net675));
 sg13g2_tiehi _08018__676 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net676));
 sg13g2_tiehi _08017__677 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net677));
 sg13g2_tiehi _08016__678 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net678));
 sg13g2_tiehi _08015__679 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net679));
 sg13g2_tiehi _08014__680 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net680));
 sg13g2_tiehi _08013__681 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net681));
 sg13g2_tiehi _08012__682 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net682));
 sg13g2_tiehi _08399__683 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net683));
 sg13g2_tiehi _08011__684 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net684));
 sg13g2_tiehi _08010__685 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net685));
 sg13g2_tiehi _08009__686 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net686));
 sg13g2_tiehi _08008__687 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net687));
 sg13g2_tiehi _08007__688 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net688));
 sg13g2_tiehi _08006__689 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net689));
 sg13g2_tiehi _08005__690 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net690));
 sg13g2_tiehi _08004__691 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net691));
 sg13g2_tiehi _08003__692 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net692));
 sg13g2_tiehi _08002__693 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net693));
 sg13g2_tiehi _08001__694 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net694));
 sg13g2_tiehi _08000__695 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net695));
 sg13g2_tiehi _07999__696 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net696));
 sg13g2_tiehi _09239__697 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net697));
 sg13g2_tiehi _07958__698 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net698));
 sg13g2_tiehi _09238__699 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net699));
 sg13g2_tiehi _07957__700 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net700));
 sg13g2_tiehi _09237__701 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net701));
 sg13g2_tiehi _08553__702 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net702));
 sg13g2_tiehi _07956__703 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net703));
 sg13g2_tiehi _09236__704 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net704));
 sg13g2_tiehi _07955__705 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net705));
 sg13g2_tiehi _07950__706 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net706));
 sg13g2_tiehi _07949__707 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net707));
 sg13g2_tiehi _07948__708 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net708));
 sg13g2_tiehi _07939__709 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net709));
 sg13g2_tiehi _07938__710 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net710));
 sg13g2_tiehi _07937__711 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net711));
 sg13g2_tiehi _07936__712 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net712));
 sg13g2_tiehi _07935__713 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net713));
 sg13g2_tiehi _07934__714 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net714));
 sg13g2_tiehi _07933__715 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net715));
 sg13g2_tiehi _07932__716 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net716));
 sg13g2_tiehi _07931__717 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net717));
 sg13g2_tiehi _07930__718 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net718));
 sg13g2_tiehi _07929__719 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net719));
 sg13g2_tiehi _07928__720 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net720));
 sg13g2_tiehi _07927__721 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net721));
 sg13g2_tiehi _07926__722 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net722));
 sg13g2_tiehi _07925__723 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net723));
 sg13g2_tiehi _07924__724 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net724));
 sg13g2_tiehi _07923__725 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net725));
 sg13g2_tiehi _07922__726 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net726));
 sg13g2_tiehi _07921__727 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net727));
 sg13g2_tiehi _07920__728 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net728));
 sg13g2_tiehi _07919__729 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net729));
 sg13g2_tiehi _07918__730 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net730));
 sg13g2_tiehi _07917__731 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net731));
 sg13g2_tiehi _07916__732 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net732));
 sg13g2_tiehi _07915__733 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net733));
 sg13g2_tiehi _07914__734 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net734));
 sg13g2_tiehi _07913__735 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net735));
 sg13g2_tiehi _07912__736 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net736));
 sg13g2_tiehi _07911__737 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net737));
 sg13g2_tiehi _07910__738 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net738));
 sg13g2_tiehi _07909__739 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net739));
 sg13g2_tiehi _08586__740 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net740));
 sg13g2_tiehi _08626__741 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net741));
 sg13g2_tiehi _08627__742 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net742));
 sg13g2_tiehi _08628__743 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net743));
 sg13g2_tiehi _09235__744 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net744));
 sg13g2_tiehi _09234__745 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net745));
 sg13g2_tiehi _09233__746 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net746));
 sg13g2_tiehi _09232__747 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net747));
 sg13g2_tiehi _09231__748 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net748));
 sg13g2_tiehi _09230__749 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net749));
 sg13g2_tiehi _09229__750 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net750));
 sg13g2_tiehi _09228__751 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net751));
 sg13g2_tiehi _09227__752 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net752));
 sg13g2_tiehi _09226__753 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net753));
 sg13g2_tiehi _09225__754 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net754));
 sg13g2_tiehi _09224__755 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net755));
 sg13g2_tiehi _09223__756 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net756));
 sg13g2_tiehi _09222__757 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net757));
 sg13g2_tiehi _09221__758 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net758));
 sg13g2_tiehi _09220__759 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net759));
 sg13g2_tiehi _09219__760 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net760));
 sg13g2_tiehi _09218__761 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net761));
 sg13g2_tiehi _09217__762 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net762));
 sg13g2_tiehi _09216__763 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net763));
 sg13g2_tiehi _09215__764 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net764));
 sg13g2_tiehi _09214__765 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net765));
 sg13g2_tiehi _09213__766 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net766));
 sg13g2_tiehi _09212__767 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net767));
 sg13g2_tiehi _09211__768 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net768));
 sg13g2_tiehi _09210__769 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net769));
 sg13g2_tiehi _09209__770 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net770));
 sg13g2_tiehi _09208__771 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net771));
 sg13g2_tiehi _09207__772 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net772));
 sg13g2_tiehi _09206__773 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net773));
 sg13g2_tiehi _08629__774 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net774));
 sg13g2_tiehi _08662__775 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net775));
 sg13g2_tiehi _09205__776 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net776));
 sg13g2_tiehi _09204__777 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net777));
 sg13g2_tiehi _09203__778 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net778));
 sg13g2_tiehi _09202__779 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net779));
 sg13g2_tiehi _09201__780 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net780));
 sg13g2_tiehi _09200__781 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net781));
 sg13g2_tiehi _09199__782 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net782));
 sg13g2_tiehi _09198__783 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net783));
 sg13g2_tiehi _09197__784 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net784));
 sg13g2_tiehi _09196__785 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net785));
 sg13g2_tiehi _09195__786 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net786));
 sg13g2_tiehi _09194__787 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net787));
 sg13g2_tiehi _09193__788 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net788));
 sg13g2_tiehi _09192__789 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net789));
 sg13g2_tiehi _09191__790 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net790));
 sg13g2_tiehi _09190__791 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net791));
 sg13g2_tiehi _09189__792 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net792));
 sg13g2_tiehi _09188__793 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net793));
 sg13g2_tiehi _09187__794 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net794));
 sg13g2_tiehi _09186__795 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net795));
 sg13g2_tiehi _09185__796 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net796));
 sg13g2_tiehi _09184__797 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net797));
 sg13g2_tiehi _09183__798 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net798));
 sg13g2_tiehi _09182__799 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net799));
 sg13g2_tiehi _09181__800 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net800));
 sg13g2_tiehi _09180__801 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net801));
 sg13g2_tiehi _09179__802 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net802));
 sg13g2_tiehi _09178__803 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net803));
 sg13g2_tiehi _09048__804 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net804));
 sg13g2_tiehi _09177__805 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net805));
 sg13g2_tiehi _09176__806 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net806));
 sg13g2_tiehi _09175__807 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net807));
 sg13g2_tiehi _09174__808 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net808));
 sg13g2_tiehi _09173__809 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net809));
 sg13g2_tiehi _09172__810 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net810));
 sg13g2_tiehi _09171__811 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net811));
 sg13g2_tiehi _09170__812 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net812));
 sg13g2_tiehi _09169__813 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net813));
 sg13g2_tiehi _09168__814 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net814));
 sg13g2_tiehi _09167__815 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net815));
 sg13g2_tiehi _09166__816 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net816));
 sg13g2_tiehi _09165__817 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net817));
 sg13g2_tiehi _09164__818 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net818));
 sg13g2_tiehi _09163__819 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net819));
 sg13g2_tiehi _09162__820 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net820));
 sg13g2_tiehi _09161__821 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net821));
 sg13g2_tiehi _09160__822 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net822));
 sg13g2_tiehi _09159__823 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net823));
 sg13g2_tiehi _09158__824 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net824));
 sg13g2_tiehi _09157__825 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net825));
 sg13g2_tiehi _09156__826 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net826));
 sg13g2_tiehi _09155__827 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net827));
 sg13g2_tiehi _09154__828 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net828));
 sg13g2_tiehi _09153__829 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net829));
 sg13g2_tiehi _09152__830 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net830));
 sg13g2_tiehi _09151__831 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net831));
 sg13g2_tiehi _09150__832 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net832));
 sg13g2_tiehi _09149__833 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net833));
 sg13g2_tiehi _09148__834 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net834));
 sg13g2_tiehi _09147__835 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net835));
 sg13g2_tiehi _09146__836 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net836));
 sg13g2_tiehi _09145__837 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net837));
 sg13g2_tiehi _09144__838 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net838));
 sg13g2_tiehi _09143__839 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net839));
 sg13g2_tiehi _09142__840 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net840));
 sg13g2_tiehi _09141__841 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net841));
 sg13g2_tiehi _09140__842 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net842));
 sg13g2_tiehi _09139__843 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net843));
 sg13g2_tiehi _09138__844 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net844));
 sg13g2_tiehi _09137__845 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net845));
 sg13g2_tiehi _09136__846 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net846));
 sg13g2_tiehi _09135__847 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net847));
 sg13g2_tiehi _09134__848 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net848));
 sg13g2_tiehi _09133__849 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net849));
 sg13g2_tiehi _09132__850 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net850));
 sg13g2_tiehi _09131__851 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net851));
 sg13g2_tiehi _09130__852 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net852));
 sg13g2_tiehi _09129__853 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net853));
 sg13g2_tiehi _09128__854 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net854));
 sg13g2_tiehi _09127__855 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net855));
 sg13g2_tiehi _09126__856 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net856));
 sg13g2_tiehi _09125__857 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net857));
 sg13g2_tiehi _09124__858 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net858));
 sg13g2_tiehi _09123__859 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net859));
 sg13g2_tiehi _09122__860 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net860));
 sg13g2_tiehi _09121__861 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net861));
 sg13g2_tiehi _09120__862 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net862));
 sg13g2_tiehi _09119__863 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net863));
 sg13g2_tiehi _09118__864 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net864));
 sg13g2_tiehi _09117__865 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net865));
 sg13g2_tiehi _09116__866 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net866));
 sg13g2_tiehi _09115__867 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net867));
 sg13g2_tiehi _09114__868 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net868));
 sg13g2_tiehi _09113__869 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net869));
 sg13g2_tiehi _09112__870 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net870));
 sg13g2_tiehi _09111__871 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net871));
 sg13g2_tiehi _09110__872 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1292));
 sg13g2_tiehi _09109__873 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1293));
 sg13g2_tiehi _09108__874 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1294));
 sg13g2_tiehi _09107__875 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1295));
 sg13g2_tiehi _09106__876 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1296));
 sg13g2_tiehi _09105__877 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1297));
 sg13g2_tiehi _09104__878 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1298));
 sg13g2_tiehi _09103__879 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1299));
 sg13g2_tiehi _09102__880 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1300));
 sg13g2_tiehi _09101__881 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1301));
 sg13g2_tiehi _09100__882 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1302));
 sg13g2_tiehi _09099__883 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1303));
 sg13g2_tiehi _09098__884 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1304));
 sg13g2_tiehi _09097__885 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1305));
 sg13g2_tiehi _09096__886 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1306));
 sg13g2_tiehi _09095__887 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1307));
 sg13g2_tiehi _09094__888 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1308));
 sg13g2_tiehi _09093__889 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1309));
 sg13g2_tiehi _09092__890 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1310));
 sg13g2_tiehi _09091__891 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1311));
 sg13g2_tiehi _09090__892 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1312));
 sg13g2_tiehi _09089__893 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1313));
 sg13g2_tiehi _09088__894 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1314));
 sg13g2_tiehi _09087__895 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1315));
 sg13g2_tiehi _09086__896 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1316));
 sg13g2_tiehi _09085__897 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1317));
 sg13g2_tiehi _09084__898 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1318));
 sg13g2_tiehi _09083__899 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1319));
 sg13g2_tiehi _09082__900 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1320));
 sg13g2_tiehi _09081__901 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1321));
 sg13g2_tiehi _09080__902 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1322));
 sg13g2_tiehi _09079__903 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1323));
 sg13g2_tiehi _09078__904 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1324));
 sg13g2_tiehi _09077__905 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1325));
 sg13g2_tiehi _09076__906 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1326));
 sg13g2_tiehi _09075__907 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1327));
 sg13g2_tiehi _09074__908 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1328));
 sg13g2_tiehi _09073__909 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1329));
 sg13g2_tiehi _09072__910 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1330));
 sg13g2_tiehi _09071__911 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1331));
 sg13g2_tiehi _09070__912 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1332));
 sg13g2_tiehi _09069__913 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1333));
 sg13g2_tiehi _09068__914 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1334));
 sg13g2_tiehi _09067__915 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1335));
 sg13g2_tiehi _09066__916 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1336));
 sg13g2_tiehi _09065__917 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1337));
 sg13g2_tiehi _09064__918 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1338));
 sg13g2_tiehi _09063__919 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1339));
 sg13g2_tiehi _09062__920 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1340));
 sg13g2_tiehi _09061__921 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1341));
 sg13g2_tiehi _09060__922 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1342));
 sg13g2_tiehi _09059__923 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1343));
 sg13g2_tiehi _09058__924 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1344));
 sg13g2_tiehi _09057__925 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1345));
 sg13g2_tiehi _09056__926 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1346));
 sg13g2_tiehi _09055__927 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1347));
 sg13g2_tiehi _09054__928 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1348));
 sg13g2_tiehi _09053__929 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1349));
 sg13g2_tiehi _09052__930 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1350));
 sg13g2_tiehi _09051__931 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1351));
 sg13g2_tiehi _09050__932 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1352));
 sg13g2_tiehi _09305__933 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1353));
 sg13g2_tiehi _09049__934 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1354));
 sg13g2_tiehi _09304__935 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1355));
 sg13g2_tiehi _09046__936 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1356));
 sg13g2_tiehi _09303__937 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1357));
 sg13g2_tiehi _09045__938 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1358));
 sg13g2_tiehi _09044__939 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1359));
 sg13g2_tiehi _09042__940 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1360));
 sg13g2_tiehi _09041__941 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1361));
 sg13g2_tiehi _09040__942 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1362));
 sg13g2_tiehi _09039__943 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1363));
 sg13g2_tiehi _09038__944 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1364));
 sg13g2_tiehi _09037__945 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1365));
 sg13g2_tiehi _09036__946 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1366));
 sg13g2_tiehi _09035__947 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1367));
 sg13g2_tiehi _09034__948 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1368));
 sg13g2_tiehi _09033__949 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1369));
 sg13g2_tiehi _09032__950 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1370));
 sg13g2_tiehi _09031__951 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1371));
 sg13g2_tiehi _09030__952 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1372));
 sg13g2_tiehi _09029__953 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1373));
 sg13g2_tiehi _09028__954 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1374));
 sg13g2_tiehi _09027__955 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1375));
 sg13g2_tiehi _09026__956 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1376));
 sg13g2_tiehi _09025__957 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1377));
 sg13g2_tiehi _09024__958 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1378));
 sg13g2_tiehi _09023__959 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1379));
 sg13g2_tiehi _09022__960 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1380));
 sg13g2_tiehi _09021__961 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1381));
 sg13g2_tiehi _09020__962 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1382));
 sg13g2_tiehi _09019__963 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1383));
 sg13g2_tiehi _09018__964 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1384));
 sg13g2_tiehi _09017__965 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1385));
 sg13g2_tiehi _09016__966 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1386));
 sg13g2_tiehi _09015__967 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1387));
 sg13g2_tiehi _09014__968 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1388));
 sg13g2_tiehi _09013__969 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1389));
 sg13g2_tiehi _09012__970 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1390));
 sg13g2_tiehi _09011__971 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1391));
 sg13g2_tiehi _09010__972 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1392));
 sg13g2_tiehi _09009__973 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1393));
 sg13g2_tiehi _09008__974 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1394));
 sg13g2_tiehi _09007__975 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1395));
 sg13g2_tiehi _09006__976 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1396));
 sg13g2_tiehi _09005__977 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1397));
 sg13g2_tiehi _09004__978 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1398));
 sg13g2_tiehi _09003__979 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1399));
 sg13g2_tiehi _09002__980 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1400));
 sg13g2_tiehi _09001__981 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1401));
 sg13g2_tiehi _09000__982 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1402));
 sg13g2_tiehi _08999__983 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1403));
 sg13g2_tiehi _08998__984 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1404));
 sg13g2_tiehi _08997__985 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1405));
 sg13g2_tiehi _08996__986 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1406));
 sg13g2_tiehi _08995__987 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1407));
 sg13g2_tiehi _08994__988 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1408));
 sg13g2_tiehi _08993__989 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1409));
 sg13g2_tiehi _08992__990 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1410));
 sg13g2_tiehi _08991__991 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1411));
 sg13g2_tiehi _08990__992 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1412));
 sg13g2_tiehi _08989__993 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1413));
 sg13g2_tiehi _08988__994 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1414));
 sg13g2_tiehi _08987__995 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1415));
 sg13g2_tiehi _08986__996 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1416));
 sg13g2_tiehi _08985__997 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1417));
 sg13g2_tiehi _08984__998 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1418));
 sg13g2_tiehi _08983__999 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1419));
 sg13g2_tiehi _08982__1000 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1420));
 sg13g2_tiehi _08981__1001 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1421));
 sg13g2_tiehi _08980__1002 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1422));
 sg13g2_tiehi _08979__1003 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1423));
 sg13g2_tiehi _08978__1004 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1424));
 sg13g2_tiehi _08977__1005 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1425));
 sg13g2_tiehi _08976__1006 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1426));
 sg13g2_tiehi _08975__1007 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1427));
 sg13g2_tiehi _08974__1008 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1428));
 sg13g2_tiehi _08973__1009 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1429));
 sg13g2_tiehi _08972__1010 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1430));
 sg13g2_tiehi _08971__1011 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1431));
 sg13g2_tiehi _08970__1012 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1432));
 sg13g2_tiehi _08969__1013 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1433));
 sg13g2_tiehi _08968__1014 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1434));
 sg13g2_tiehi _08967__1015 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1435));
 sg13g2_tiehi _08966__1016 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1436));
 sg13g2_tiehi _08965__1017 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1437));
 sg13g2_tiehi _08964__1018 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1438));
 sg13g2_tiehi _08963__1019 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1439));
 sg13g2_tiehi _08962__1020 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1440));
 sg13g2_tiehi _08961__1021 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1441));
 sg13g2_tiehi _08960__1022 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1442));
 sg13g2_tiehi _08959__1023 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1443));
 sg13g2_tiehi _08958__1024 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1444));
 sg13g2_tiehi _08957__1025 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1445));
 sg13g2_tiehi _08956__1026 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1446));
 sg13g2_tiehi _08955__1027 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1447));
 sg13g2_tiehi _08954__1028 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1448));
 sg13g2_tiehi _08953__1029 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1449));
 sg13g2_tiehi _08952__1030 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1450));
 sg13g2_tiehi _08951__1031 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1451));
 sg13g2_tiehi _08950__1032 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1452));
 sg13g2_tiehi _08949__1033 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1453));
 sg13g2_tiehi _08948__1034 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1454));
 sg13g2_tiehi _08947__1035 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1455));
 sg13g2_tiehi _08946__1036 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1456));
 sg13g2_tiehi _08945__1037 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1457));
 sg13g2_tiehi _08944__1038 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1458));
 sg13g2_tiehi _08943__1039 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1459));
 sg13g2_tiehi _08942__1040 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1460));
 sg13g2_tiehi _08941__1041 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1461));
 sg13g2_tiehi _08940__1042 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1462));
 sg13g2_tiehi _08939__1043 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1463));
 sg13g2_tiehi _08938__1044 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1464));
 sg13g2_tiehi _08937__1045 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1465));
 sg13g2_tiehi _08936__1046 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1466));
 sg13g2_tiehi _08935__1047 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1467));
 sg13g2_tiehi _08934__1048 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1468));
 sg13g2_tiehi _08933__1049 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1469));
 sg13g2_tiehi _08932__1050 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1470));
 sg13g2_tiehi _08931__1051 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1471));
 sg13g2_tiehi _08930__1052 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1472));
 sg13g2_tiehi _08929__1053 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1473));
 sg13g2_tiehi _08928__1054 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1474));
 sg13g2_tiehi _08927__1055 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1475));
 sg13g2_tiehi _08926__1056 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1476));
 sg13g2_tiehi _08925__1057 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1477));
 sg13g2_tiehi _08924__1058 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1478));
 sg13g2_tiehi _08923__1059 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1479));
 sg13g2_tiehi _08922__1060 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1480));
 sg13g2_tiehi _08921__1061 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1481));
 sg13g2_tiehi _08920__1062 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1482));
 sg13g2_tiehi _08919__1063 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1483));
 sg13g2_tiehi _08918__1064 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1484));
 sg13g2_tiehi _08917__1065 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1485));
 sg13g2_tiehi _08916__1066 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1486));
 sg13g2_tiehi _08915__1067 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1487));
 sg13g2_tiehi _08914__1068 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1488));
 sg13g2_tiehi _08913__1069 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1489));
 sg13g2_tiehi _08912__1070 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1490));
 sg13g2_tiehi _08911__1071 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1491));
 sg13g2_tiehi _08910__1072 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1492));
 sg13g2_tiehi _08909__1073 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1493));
 sg13g2_tiehi _08908__1074 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1494));
 sg13g2_tiehi _08907__1075 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1495));
 sg13g2_tiehi _08906__1076 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1496));
 sg13g2_tiehi _08905__1077 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1497));
 sg13g2_tiehi _08904__1078 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1498));
 sg13g2_tiehi _08903__1079 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1499));
 sg13g2_tiehi _08902__1080 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1500));
 sg13g2_tiehi _08901__1081 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1501));
 sg13g2_tiehi _08900__1082 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1502));
 sg13g2_tiehi _08899__1083 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1503));
 sg13g2_tiehi _08898__1084 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1504));
 sg13g2_tiehi _08897__1085 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1505));
 sg13g2_tiehi _08896__1086 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1506));
 sg13g2_tiehi _08895__1087 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1507));
 sg13g2_tiehi _08894__1088 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1508));
 sg13g2_tiehi _08893__1089 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1509));
 sg13g2_tiehi _08892__1090 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1510));
 sg13g2_tiehi _08891__1091 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1511));
 sg13g2_tiehi _08890__1092 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1512));
 sg13g2_tiehi _08889__1093 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1513));
 sg13g2_tiehi _08888__1094 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1514));
 sg13g2_tiehi _08887__1095 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1515));
 sg13g2_tiehi _08886__1096 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1516));
 sg13g2_tiehi _08885__1097 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1517));
 sg13g2_tiehi _08884__1098 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1518));
 sg13g2_tiehi _08883__1099 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1519));
 sg13g2_tiehi _08882__1100 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1520));
 sg13g2_tiehi _08881__1101 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1521));
 sg13g2_tiehi _08880__1102 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1522));
 sg13g2_tiehi _08879__1103 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1523));
 sg13g2_tiehi _08878__1104 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1524));
 sg13g2_tiehi _08877__1105 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1525));
 sg13g2_tiehi _08876__1106 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1526));
 sg13g2_tiehi _08875__1107 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1527));
 sg13g2_tiehi _08874__1108 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1528));
 sg13g2_tiehi _08873__1109 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1529));
 sg13g2_tiehi _08872__1110 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1530));
 sg13g2_tiehi _08871__1111 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1531));
 sg13g2_tiehi _08870__1112 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1532));
 sg13g2_tiehi _09302__1113 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1533));
 sg13g2_tiehi _08869__1114 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1534));
 sg13g2_tiehi _09301__1115 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1535));
 sg13g2_tiehi _08868__1116 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1536));
 sg13g2_tiehi _09300__1117 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1537));
 sg13g2_tiehi _08867__1118 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1538));
 sg13g2_tiehi _09299__1119 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1539));
 sg13g2_tiehi _08866__1120 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1540));
 sg13g2_tiehi _08865__1121 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1541));
 sg13g2_tiehi _08864__1122 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1542));
 sg13g2_tiehi _08863__1123 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1543));
 sg13g2_tiehi _08862__1124 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1544));
 sg13g2_tiehi _08861__1125 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1545));
 sg13g2_tiehi _08860__1126 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1546));
 sg13g2_tiehi _08859__1127 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1547));
 sg13g2_tiehi _08858__1128 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1548));
 sg13g2_tiehi _08857__1129 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1549));
 sg13g2_tiehi _08856__1130 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1550));
 sg13g2_tiehi _08855__1131 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1551));
 sg13g2_tiehi _08854__1132 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1552));
 sg13g2_tiehi _08853__1133 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1553));
 sg13g2_tiehi _08852__1134 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1554));
 sg13g2_tiehi _08851__1135 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1555));
 sg13g2_tiehi _08850__1136 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1556));
 sg13g2_tiehi _08849__1137 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1557));
 sg13g2_tiehi _08848__1138 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1558));
 sg13g2_tiehi _08847__1139 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1559));
 sg13g2_tiehi _08846__1140 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1560));
 sg13g2_tiehi _08845__1141 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1561));
 sg13g2_tiehi _08844__1142 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1562));
 sg13g2_tiehi _08843__1143 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1563));
 sg13g2_tiehi _08842__1144 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1564));
 sg13g2_tiehi _08841__1145 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1565));
 sg13g2_tiehi _08840__1146 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1566));
 sg13g2_tiehi _08839__1147 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1567));
 sg13g2_tiehi _08838__1148 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1568));
 sg13g2_tiehi _08837__1149 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1569));
 sg13g2_tiehi _09043__1150 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1570));
 sg13g2_tiehi _09047__1151 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1571));
 sg13g2_tiehi _08836__1152 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1572));
 sg13g2_tiehi _08835__1153 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1573));
 sg13g2_tiehi _08834__1154 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1574));
 sg13g2_tiehi _08833__1155 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1575));
 sg13g2_tiehi _08832__1156 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1576));
 sg13g2_tiehi _08831__1157 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1577));
 sg13g2_tiehi _08830__1158 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1578));
 sg13g2_tiehi _08829__1159 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1579));
 sg13g2_tiehi _08828__1160 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1580));
 sg13g2_tiehi _08827__1161 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1581));
 sg13g2_tiehi _08826__1162 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1582));
 sg13g2_tiehi _08825__1163 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1583));
 sg13g2_tiehi _08824__1164 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1584));
 sg13g2_tiehi _08823__1165 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1585));
 sg13g2_tiehi _08822__1166 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1586));
 sg13g2_tiehi _08821__1167 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1587));
 sg13g2_tiehi _08820__1168 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1588));
 sg13g2_tiehi _08819__1169 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1589));
 sg13g2_tiehi _08818__1170 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1590));
 sg13g2_tiehi _08817__1171 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1591));
 sg13g2_tiehi _08816__1172 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1592));
 sg13g2_tiehi _08815__1173 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1593));
 sg13g2_tiehi _08814__1174 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1594));
 sg13g2_tiehi _08813__1175 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1595));
 sg13g2_tiehi _08812__1176 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1596));
 sg13g2_tiehi _08811__1177 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1597));
 sg13g2_tiehi _08810__1178 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1598));
 sg13g2_tiehi _08809__1179 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1599));
 sg13g2_tiehi _08808__1180 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1600));
 sg13g2_tiehi _08807__1181 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1601));
 sg13g2_tiehi _08806__1182 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1602));
 sg13g2_tiehi _08805__1183 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1603));
 sg13g2_tiehi _08804__1184 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1604));
 sg13g2_tiehi _08803__1185 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1605));
 sg13g2_tiehi _08802__1186 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1606));
 sg13g2_tiehi _08801__1187 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1607));
 sg13g2_tiehi _08800__1188 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1608));
 sg13g2_tiehi _08799__1189 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1609));
 sg13g2_tiehi _08798__1190 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1610));
 sg13g2_tiehi _08797__1191 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1611));
 sg13g2_tiehi _08796__1192 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1612));
 sg13g2_tiehi _08795__1193 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1613));
 sg13g2_tiehi _08794__1194 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1614));
 sg13g2_tiehi _08793__1195 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1615));
 sg13g2_tiehi _08792__1196 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1616));
 sg13g2_tiehi _08791__1197 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1617));
 sg13g2_tiehi _08790__1198 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1618));
 sg13g2_tiehi _08789__1199 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1619));
 sg13g2_tiehi _08788__1200 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1620));
 sg13g2_tiehi _08787__1201 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1621));
 sg13g2_tiehi _08786__1202 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1622));
 sg13g2_tiehi _08785__1203 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1623));
 sg13g2_tiehi _08784__1204 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1624));
 sg13g2_tiehi _08783__1205 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1625));
 sg13g2_tiehi _08782__1206 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1626));
 sg13g2_tiehi _08781__1207 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1627));
 sg13g2_tiehi _08780__1208 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1628));
 sg13g2_tiehi _08779__1209 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1629));
 sg13g2_tiehi _08778__1210 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1630));
 sg13g2_tiehi _08777__1211 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1631));
 sg13g2_tiehi _08776__1212 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1632));
 sg13g2_tiehi _08775__1213 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1633));
 sg13g2_tiehi _08774__1214 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1634));
 sg13g2_tiehi _08773__1215 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1635));
 sg13g2_tiehi _08772__1216 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1636));
 sg13g2_tiehi _08771__1217 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1637));
 sg13g2_tiehi _08770__1218 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1638));
 sg13g2_tiehi _08769__1219 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1639));
 sg13g2_tiehi _08768__1220 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1640));
 sg13g2_tiehi _08767__1221 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1641));
 sg13g2_tiehi _08766__1222 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1642));
 sg13g2_tiehi _08765__1223 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1643));
 sg13g2_tiehi _08764__1224 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1644));
 sg13g2_tiehi _08763__1225 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1645));
 sg13g2_tiehi _08762__1226 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1646));
 sg13g2_tiehi _08761__1227 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1647));
 sg13g2_tiehi _08760__1228 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1648));
 sg13g2_tiehi _08759__1229 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1649));
 sg13g2_tiehi _08758__1230 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1650));
 sg13g2_tiehi _08757__1231 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1651));
 sg13g2_tiehi _08756__1232 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1652));
 sg13g2_tiehi _08755__1233 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1653));
 sg13g2_tiehi _08754__1234 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1654));
 sg13g2_tiehi _08753__1235 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1655));
 sg13g2_tiehi _08752__1236 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1656));
 sg13g2_tiehi _08751__1237 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1657));
 sg13g2_tiehi _08750__1238 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1658));
 sg13g2_tiehi _08749__1239 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1659));
 sg13g2_tiehi _08748__1240 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1660));
 sg13g2_tiehi _08747__1241 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1661));
 sg13g2_tiehi _08746__1242 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1662));
 sg13g2_tiehi _08745__1243 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1663));
 sg13g2_tiehi _08744__1244 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1664));
 sg13g2_tiehi _08743__1245 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1665));
 sg13g2_tiehi _08742__1246 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1666));
 sg13g2_tiehi _08741__1247 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1667));
 sg13g2_tiehi _08740__1248 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1668));
 sg13g2_tiehi _08739__1249 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1669));
 sg13g2_tiehi _08738__1250 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1670));
 sg13g2_tiehi _08737__1251 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1671));
 sg13g2_tiehi _08736__1252 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1672));
 sg13g2_tiehi _08735__1253 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1673));
 sg13g2_tiehi _08734__1254 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1674));
 sg13g2_tiehi _08733__1255 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1675));
 sg13g2_tiehi _08732__1256 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1676));
 sg13g2_tiehi _08731__1257 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1677));
 sg13g2_tiehi _08730__1258 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1678));
 sg13g2_tiehi _08729__1259 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1679));
 sg13g2_tiehi _08728__1260 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1680));
 sg13g2_tiehi _08727__1261 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1681));
 sg13g2_tiehi _08726__1262 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1682));
 sg13g2_tiehi _08725__1263 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1683));
 sg13g2_tiehi _08724__1264 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1684));
 sg13g2_tiehi _08723__1265 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1685));
 sg13g2_tiehi _08722__1266 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1686));
 sg13g2_tiehi _08721__1267 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1687));
 sg13g2_tiehi _08720__1268 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1688));
 sg13g2_tiehi _08719__1269 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1689));
 sg13g2_tiehi _08718__1270 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1690));
 sg13g2_tiehi _08717__1271 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1691));
 sg13g2_tiehi _08716__1272 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1692));
 sg13g2_tiehi _08715__1273 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1693));
 sg13g2_tiehi _08714__1274 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1694));
 sg13g2_tiehi _08713__1275 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1695));
 sg13g2_tiehi _08712__1276 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1696));
 sg13g2_tiehi _08711__1277 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1697));
 sg13g2_tiehi _08710__1278 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1698));
 sg13g2_tiehi _08709__1279 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1699));
 sg13g2_tiehi _08708__1280 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1700));
 sg13g2_tiehi _08707__1281 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1701));
 sg13g2_tiehi _08706__1282 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1702));
 sg13g2_tiehi _08705__1283 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1703));
 sg13g2_tiehi _08704__1284 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1704));
 sg13g2_tiehi _08703__1285 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1705));
 sg13g2_tiehi _08702__1286 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1706));
 sg13g2_tiehi _08701__1287 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1707));
 sg13g2_tiehi _08700__1288 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1708));
 sg13g2_tiehi _08699__1289 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1709));
 sg13g2_tiehi _08698__1290 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1710));
 sg13g2_tiehi _08697__1291 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1711));
 sg13g2_tiehi _08696__1292 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1712));
 sg13g2_tiehi _08695__1293 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1713));
 sg13g2_tiehi _08694__1294 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1714));
 sg13g2_tiehi _08693__1295 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1715));
 sg13g2_tiehi _08692__1296 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1716));
 sg13g2_tiehi _08691__1297 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1717));
 sg13g2_tiehi _08690__1298 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1718));
 sg13g2_tiehi _08689__1299 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1719));
 sg13g2_tiehi _08688__1300 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1720));
 sg13g2_tiehi _08687__1301 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1721));
 sg13g2_tiehi _08686__1302 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1722));
 sg13g2_tiehi _08685__1303 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1723));
 sg13g2_tiehi _08684__1304 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1724));
 sg13g2_tiehi _08683__1305 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1725));
 sg13g2_tiehi _08682__1306 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1726));
 sg13g2_tiehi _08681__1307 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1727));
 sg13g2_tiehi _08680__1308 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1728));
 sg13g2_tiehi _08679__1309 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1729));
 sg13g2_tiehi _08678__1310 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1730));
 sg13g2_tiehi _08677__1311 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1731));
 sg13g2_tiehi _08676__1312 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1732));
 sg13g2_tiehi _08675__1313 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1733));
 sg13g2_tiehi _08674__1314 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1734));
 sg13g2_tiehi _08673__1315 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1735));
 sg13g2_tiehi _08661__1316 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1736));
 sg13g2_tiehi _08660__1317 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1737));
 sg13g2_tiehi _08659__1318 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1738));
 sg13g2_tiehi _08658__1319 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1739));
 sg13g2_tiehi _08657__1320 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1740));
 sg13g2_tiehi _08656__1321 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1741));
 sg13g2_tiehi _08655__1322 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1742));
 sg13g2_tiehi _08654__1323 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1743));
 sg13g2_tiehi _08653__1324 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1744));
 sg13g2_tiehi _08652__1325 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1745));
 sg13g2_tiehi _08651__1326 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1746));
 sg13g2_tiehi _08650__1327 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1747));
 sg13g2_tiehi _08649__1328 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1748));
 sg13g2_tiehi _08648__1329 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1749));
 sg13g2_tiehi _08647__1330 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1750));
 sg13g2_tiehi _08646__1331 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1751));
 sg13g2_tiehi _08645__1332 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1752));
 sg13g2_tiehi _08644__1333 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1753));
 sg13g2_tiehi _08643__1334 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1754));
 sg13g2_tiehi _08642__1335 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1755));
 sg13g2_tiehi _08641__1336 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1756));
 sg13g2_tiehi _08640__1337 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1757));
 sg13g2_tiehi _08639__1338 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1758));
 sg13g2_tiehi _08638__1339 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1759));
 sg13g2_tiehi _08637__1340 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1760));
 sg13g2_tiehi _08636__1341 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1761));
 sg13g2_tiehi _08635__1342 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1762));
 sg13g2_tiehi _08634__1343 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1763));
 sg13g2_tiehi _08633__1344 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1764));
 sg13g2_tiehi _08632__1345 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1765));
 sg13g2_tiehi _08631__1346 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1766));
 sg13g2_tiehi _09298__1347 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1767));
 sg13g2_tiehi _08630__1348 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1768));
 sg13g2_tiehi _09297__1349 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1769));
 sg13g2_tiehi _08625__1350 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1770));
 sg13g2_tiehi _09296__1351 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1771));
 sg13g2_tiehi _08624__1352 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1772));
 sg13g2_tiehi _08623__1353 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1773));
 sg13g2_tiehi _08622__1354 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1774));
 sg13g2_tiehi _08621__1355 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1775));
 sg13g2_tiehi _08620__1356 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1776));
 sg13g2_tiehi _08619__1357 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1777));
 sg13g2_tiehi _08618__1358 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1778));
 sg13g2_tiehi _08617__1359 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1779));
 sg13g2_tiehi _08616__1360 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1780));
 sg13g2_tiehi _08615__1361 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1781));
 sg13g2_tiehi _08614__1362 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1782));
 sg13g2_tiehi _08613__1363 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1783));
 sg13g2_tiehi _08612__1364 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1784));
 sg13g2_tiehi _08611__1365 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1785));
 sg13g2_tiehi _08610__1366 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1786));
 sg13g2_tiehi _08609__1367 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1787));
 sg13g2_tiehi _08608__1368 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1788));
 sg13g2_tiehi _08607__1369 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1789));
 sg13g2_tiehi _08606__1370 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1790));
 sg13g2_tiehi _08605__1371 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1791));
 sg13g2_tiehi _08604__1372 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1792));
 sg13g2_tiehi _08603__1373 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1793));
 sg13g2_tiehi _08602__1374 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1794));
 sg13g2_tiehi _08601__1375 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1795));
 sg13g2_tiehi _08600__1376 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1796));
 sg13g2_tiehi _08599__1377 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1797));
 sg13g2_tiehi _08598__1378 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1798));
 sg13g2_tiehi _08597__1379 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1799));
 sg13g2_tiehi _08596__1380 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1800));
 sg13g2_tiehi _08595__1381 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1801));
 sg13g2_tiehi _08594__1382 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1802));
 sg13g2_tiehi _08593__1383 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1803));
 sg13g2_tiehi _08592__1384 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1804));
 sg13g2_tiehi _08591__1385 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1805));
 sg13g2_tiehi _08590__1386 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1806));
 sg13g2_tiehi _08589__1387 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1807));
 sg13g2_tiehi _08588__1388 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1808));
 sg13g2_tiehi _09295__1389 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1809));
 sg13g2_tiehi _08587__1390 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1810));
 sg13g2_tiehi _09294__1391 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1811));
 sg13g2_tiehi _08585__1392 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1812));
 sg13g2_tiehi _09293__1393 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1813));
 sg13g2_tiehi _08584__1394 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1814));
 sg13g2_tiehi _09292__1395 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1815));
 sg13g2_tiehi _08583__1396 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1816));
 sg13g2_tiehi _09291__1397 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1817));
 sg13g2_tiehi _08582__1398 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1818));
 sg13g2_tiehi _09290__1399 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1819));
 sg13g2_tiehi _08581__1400 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1820));
 sg13g2_tiehi _09289__1401 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1821));
 sg13g2_tiehi _08580__1402 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1822));
 sg13g2_tiehi _09288__1403 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1823));
 sg13g2_tiehi _08579__1404 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1824));
 sg13g2_tiehi _09287__1405 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1825));
 sg13g2_tiehi _08578__1406 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net1826));
 sg13g2_inv_1 _04658__1 (.VDD(VPWR),
    .Y(net1827),
    .A(clknet_1_0__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_1 _10671_ (.A(net1246),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10672_ (.A(net22),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10673_ (.A(net22),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10674_ (.A(ccx_req),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10675_ (.A(\i_exotiny.i_wb_spi.sck_r ),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10676_ (.A(\i_exotiny.i_wb_spi.spi_sdo_o ),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10677_ (.A(\i_exotiny._5420_$func$/home/user/heichips25-fazyrv-exotiny/build/exotiny_preproc.v:7404$13.$result [0]),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10678_ (.A(net1827),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10679_ (.A(\i_exotiny._5416_$func$/home/user/heichips25-fazyrv-exotiny/build/exotiny_preproc.v:7385$12.$result [0]),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10680_ (.A(gpo),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout872 (.A(_02472_),
    .X(net872),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout873 (.A(net875),
    .X(net873),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout874 (.A(net875),
    .X(net874),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout875 (.A(_02472_),
    .X(net875),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout876 (.A(net880),
    .X(net876),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout877 (.A(net879),
    .X(net877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout878 (.A(net879),
    .X(net878),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout879 (.A(net880),
    .X(net879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout880 (.A(_02463_),
    .X(net880),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout881 (.A(net885),
    .X(net881),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout882 (.A(net884),
    .X(net882),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout883 (.A(net884),
    .X(net883),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout884 (.A(net885),
    .X(net884),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout885 (.A(_02454_),
    .X(net885),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout886 (.A(net890),
    .X(net886),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout887 (.A(net889),
    .X(net887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout888 (.A(net889),
    .X(net888),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout889 (.A(net890),
    .X(net889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout890 (.A(_02444_),
    .X(net890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout891 (.A(net892),
    .X(net891),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout892 (.A(_03217_),
    .X(net892),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout893 (.A(net895),
    .X(net893),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout894 (.A(net895),
    .X(net894),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout895 (.A(_03217_),
    .X(net895),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout896 (.A(net897),
    .X(net896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout897 (.A(net900),
    .X(net897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout898 (.A(net900),
    .X(net898),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout899 (.A(net900),
    .X(net899),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout900 (.A(_03188_),
    .X(net900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout901 (.A(net902),
    .X(net901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout902 (.A(net903),
    .X(net902),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout903 (.A(net907),
    .X(net903),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout904 (.A(net906),
    .X(net904),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout905 (.A(net906),
    .X(net905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout906 (.A(net907),
    .X(net906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout907 (.A(_03105_),
    .X(net907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout908 (.A(net912),
    .X(net908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout909 (.A(net912),
    .X(net909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout910 (.A(net912),
    .X(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout911 (.A(net912),
    .X(net911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout912 (.A(_02979_),
    .X(net912),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout913 (.A(net915),
    .X(net913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout914 (.A(net915),
    .X(net914),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout915 (.A(net917),
    .X(net915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout916 (.A(net917),
    .X(net916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout917 (.A(_02941_),
    .X(net917),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout918 (.A(net923),
    .X(net918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout919 (.A(net923),
    .X(net919),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout920 (.A(net923),
    .X(net920),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout921 (.A(net922),
    .X(net921),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout922 (.A(net923),
    .X(net922),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout923 (.A(_02929_),
    .X(net923),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout924 (.A(net928),
    .X(net924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout925 (.A(net928),
    .X(net925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout926 (.A(net928),
    .X(net926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout927 (.A(net928),
    .X(net927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout928 (.A(_02917_),
    .X(net928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout929 (.A(net931),
    .X(net929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout930 (.A(net931),
    .X(net930),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout931 (.A(_02621_),
    .X(net931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout932 (.A(_02621_),
    .X(net932),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout933 (.A(_02621_),
    .X(net933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout934 (.A(net936),
    .X(net934),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout935 (.A(net936),
    .X(net935),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout936 (.A(_02609_),
    .X(net936),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout937 (.A(net938),
    .X(net937),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout938 (.A(_02609_),
    .X(net938),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout939 (.A(net941),
    .X(net939),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout940 (.A(net941),
    .X(net940),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout941 (.A(net944),
    .X(net941),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout942 (.A(net944),
    .X(net942),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout943 (.A(net944),
    .X(net943),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout944 (.A(_02553_),
    .X(net944),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout945 (.A(net949),
    .X(net945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout946 (.A(net949),
    .X(net946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout947 (.A(net949),
    .X(net947),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout948 (.A(net949),
    .X(net948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout949 (.A(_02541_),
    .X(net949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout950 (.A(net951),
    .X(net950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout951 (.A(net954),
    .X(net951),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout952 (.A(net953),
    .X(net952),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout953 (.A(net954),
    .X(net953),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout954 (.A(_02534_),
    .X(net954),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout955 (.A(net956),
    .X(net955),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout956 (.A(net957),
    .X(net956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout957 (.A(_02520_),
    .X(net957),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout958 (.A(net959),
    .X(net958),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout959 (.A(net960),
    .X(net959),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout960 (.A(_02520_),
    .X(net960),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout961 (.A(net965),
    .X(net961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout962 (.A(net965),
    .X(net962),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout963 (.A(net964),
    .X(net963),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout964 (.A(net965),
    .X(net964),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout965 (.A(_02511_),
    .X(net965),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout966 (.A(net971),
    .X(net966),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout967 (.A(net971),
    .X(net967),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout968 (.A(net970),
    .X(net968),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout969 (.A(net971),
    .X(net969),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout970 (.A(net971),
    .X(net970),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout971 (.A(_02487_),
    .X(net971),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout972 (.A(net977),
    .X(net972),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout973 (.A(net976),
    .X(net973),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout974 (.A(net976),
    .X(net974),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout975 (.A(net976),
    .X(net975),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout976 (.A(net977),
    .X(net976),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout977 (.A(_02479_),
    .X(net977),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout978 (.A(net980),
    .X(net978),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout979 (.A(net980),
    .X(net979),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout980 (.A(_03229_),
    .X(net980),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout981 (.A(net982),
    .X(net981),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout982 (.A(_03229_),
    .X(net982),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout983 (.A(net985),
    .X(net983),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout984 (.A(net985),
    .X(net984),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout985 (.A(net987),
    .X(net985),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout986 (.A(net987),
    .X(net986),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout987 (.A(_03223_),
    .X(net987),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout988 (.A(_03211_),
    .X(net988),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout989 (.A(_03211_),
    .X(net989),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout990 (.A(net992),
    .X(net990),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout991 (.A(net992),
    .X(net991),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout992 (.A(_03211_),
    .X(net992),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout993 (.A(net994),
    .X(net993),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout994 (.A(net997),
    .X(net994),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout995 (.A(net996),
    .X(net995),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout996 (.A(net997),
    .X(net996),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout997 (.A(_03200_),
    .X(net997),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout998 (.A(net999),
    .X(net998),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout999 (.A(_03194_),
    .X(net999),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1000 (.A(net1002),
    .X(net1000),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1001 (.A(net1002),
    .X(net1001),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1002 (.A(_03194_),
    .X(net1002),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1003 (.A(net1004),
    .X(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1004 (.A(net1007),
    .X(net1004),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1005 (.A(net1006),
    .X(net1005),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1006 (.A(net1007),
    .X(net1006),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1007 (.A(_02973_),
    .X(net1007),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1008 (.A(net1009),
    .X(net1008),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1009 (.A(net1010),
    .X(net1009),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1010 (.A(_02948_),
    .X(net1010),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1011 (.A(net1012),
    .X(net1011),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1012 (.A(_02948_),
    .X(net1012),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1013 (.A(net1014),
    .X(net1013),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1014 (.A(net1016),
    .X(net1014),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1015 (.A(net1016),
    .X(net1015),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1016 (.A(_02935_),
    .X(net1016),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1017 (.A(_02935_),
    .X(net1017),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1018 (.A(net1019),
    .X(net1018),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1019 (.A(_02923_),
    .X(net1019),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1020 (.A(net1022),
    .X(net1020),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1021 (.A(_02923_),
    .X(net1021),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1022 (.A(_02923_),
    .X(net1022),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1023 (.A(net1024),
    .X(net1023),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1024 (.A(_02615_),
    .X(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1025 (.A(net1027),
    .X(net1025),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1026 (.A(net1027),
    .X(net1026),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1027 (.A(_02615_),
    .X(net1027),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1028 (.A(net1029),
    .X(net1028),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1029 (.A(net1032),
    .X(net1029),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1030 (.A(net1031),
    .X(net1030),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1031 (.A(net1032),
    .X(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1032 (.A(_02566_),
    .X(net1032),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1033 (.A(net1034),
    .X(net1033),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1034 (.A(net1037),
    .X(net1034),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1035 (.A(net1036),
    .X(net1035),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1036 (.A(net1037),
    .X(net1036),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1037 (.A(_02559_),
    .X(net1037),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1038 (.A(net1042),
    .X(net1038),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1039 (.A(net1042),
    .X(net1039),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1040 (.A(net1042),
    .X(net1040),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1041 (.A(net1042),
    .X(net1041),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1042 (.A(_02547_),
    .X(net1042),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1043 (.A(net1045),
    .X(net1043),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1044 (.A(net1045),
    .X(net1044),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1045 (.A(_02527_),
    .X(net1045),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1046 (.A(net1047),
    .X(net1046),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1047 (.A(_02527_),
    .X(net1047),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1048 (.A(net1049),
    .X(net1048),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1049 (.A(net1052),
    .X(net1049),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1050 (.A(net1052),
    .X(net1050),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1051 (.A(net1052),
    .X(net1051),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1052 (.A(_02494_),
    .X(net1052),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1053 (.A(net1055),
    .X(net1053),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1054 (.A(net1055),
    .X(net1054),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1055 (.A(_02424_),
    .X(net1055),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1056 (.A(_02424_),
    .X(net1056),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1057 (.A(_02424_),
    .X(net1057),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1058 (.A(net1059),
    .X(net1058),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1059 (.A(net1060),
    .X(net1059),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1060 (.A(net1061),
    .X(net1060),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1061 (.A(net1067),
    .X(net1061),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1062 (.A(net1063),
    .X(net1062),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1063 (.A(net1064),
    .X(net1063),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1064 (.A(net1067),
    .X(net1064),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1065 (.A(net1066),
    .X(net1065),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1066 (.A(net1067),
    .X(net1066),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1067 (.A(_02273_),
    .X(net1067),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1068 (.A(_02718_),
    .X(net1068),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1069 (.A(net1070),
    .X(net1069),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1070 (.A(_02181_),
    .X(net1070),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1071 (.A(_02181_),
    .X(net1071),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1072 (.A(_01581_),
    .X(net1072),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1073 (.A(_01581_),
    .X(net1073),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1074 (.A(net1075),
    .X(net1074),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1075 (.A(net1076),
    .X(net1075),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1076 (.A(_01526_),
    .X(net1076),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1077 (.A(_02991_),
    .X(net1077),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1078 (.A(_02991_),
    .X(net1078),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1079 (.A(net1085),
    .X(net1079),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1080 (.A(net1084),
    .X(net1080),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1081 (.A(net1084),
    .X(net1081),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1082 (.A(net1084),
    .X(net1082),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1083 (.A(net1084),
    .X(net1083),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1084 (.A(net1085),
    .X(net1084),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1085 (.A(_02990_),
    .X(net1085),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1086 (.A(net1091),
    .X(net1086),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1087 (.A(net1091),
    .X(net1087),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1088 (.A(net1090),
    .X(net1088),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1089 (.A(net1090),
    .X(net1089),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1090 (.A(net1091),
    .X(net1090),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1091 (.A(net1092),
    .X(net1091),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1092 (.A(net1093),
    .X(net1092),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1093 (.A(_02960_),
    .X(net1093),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1094 (.A(_02717_),
    .X(net1094),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1095 (.A(_02717_),
    .X(net1095),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1096 (.A(net1101),
    .X(net1096),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1097 (.A(net1099),
    .X(net1097),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1098 (.A(net1099),
    .X(net1098),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1099 (.A(net1100),
    .X(net1099),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1100 (.A(net1101),
    .X(net1100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1101 (.A(net1102),
    .X(net1101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1102 (.A(_02717_),
    .X(net1102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1103 (.A(net1104),
    .X(net1103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1104 (.A(_02502_),
    .X(net1104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1105 (.A(\i_exotiny._2160_ ),
    .X(net1105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1106 (.A(\i_exotiny._2160_ ),
    .X(net1106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1107 (.A(net1108),
    .X(net1107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1108 (.A(_01686_),
    .X(net1108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1109 (.A(_01608_),
    .X(net1109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1110 (.A(_01607_),
    .X(net1110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1111 (.A(_01577_),
    .X(net1111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1112 (.A(_02091_),
    .X(net1112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1113 (.A(_02091_),
    .X(net1113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1114 (.A(net1115),
    .X(net1114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1115 (.A(net1116),
    .X(net1115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1116 (.A(net1117),
    .X(net1116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1117 (.A(net1120),
    .X(net1117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1118 (.A(net1119),
    .X(net1118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1119 (.A(net1120),
    .X(net1119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1120 (.A(_01582_),
    .X(net1120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1121 (.A(net1122),
    .X(net1121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1122 (.A(net1123),
    .X(net1122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1123 (.A(_01582_),
    .X(net1123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1124 (.A(net1125),
    .X(net1124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1125 (.A(_01582_),
    .X(net1125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1126 (.A(_01550_),
    .X(net1126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1127 (.A(_00026_),
    .X(net1127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1128 (.A(net1136),
    .X(net1128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1129 (.A(net1136),
    .X(net1129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1130 (.A(net1131),
    .X(net1130),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1131 (.A(net1136),
    .X(net1131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1132 (.A(net1134),
    .X(net1132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1133 (.A(net1134),
    .X(net1133),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1134 (.A(net1135),
    .X(net1134),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1135 (.A(net1136),
    .X(net1135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1136 (.A(_01507_),
    .X(net1136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1137 (.A(_01507_),
    .X(net1137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1138 (.A(net1141),
    .X(net1138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1139 (.A(net1141),
    .X(net1139),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1140 (.A(net1141),
    .X(net1140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1141 (.A(net1142),
    .X(net1141),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1142 (.A(_02422_),
    .X(net1142),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1143 (.A(_02390_),
    .X(net1143),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1144 (.A(net1145),
    .X(net1144),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1145 (.A(_01549_),
    .X(net1145),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1146 (.A(_01484_),
    .X(net1146),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1147 (.A(_03050_),
    .X(net1147),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1148 (.A(_03014_),
    .X(net1148),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1149 (.A(_03014_),
    .X(net1149),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1150 (.A(net1151),
    .X(net1150),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1151 (.A(_02984_),
    .X(net1151),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1152 (.A(net1153),
    .X(net1152),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1153 (.A(net1154),
    .X(net1153),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1154 (.A(net1157),
    .X(net1154),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1155 (.A(net1156),
    .X(net1155),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1156 (.A(net1157),
    .X(net1156),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1157 (.A(net1158),
    .X(net1157),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1158 (.A(_02415_),
    .X(net1158),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1159 (.A(net1160),
    .X(net1159),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1160 (.A(net1162),
    .X(net1160),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1161 (.A(net1162),
    .X(net1161),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1162 (.A(net1164),
    .X(net1162),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1163 (.A(net1164),
    .X(net1163),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1164 (.A(_02414_),
    .X(net1164),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1165 (.A(net1168),
    .X(net1165),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1166 (.A(net1168),
    .X(net1166),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1167 (.A(net1168),
    .X(net1167),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1168 (.A(_02414_),
    .X(net1168),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1169 (.A(_01517_),
    .X(net1169),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1170 (.A(net1171),
    .X(net1170),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1171 (.A(net1172),
    .X(net1171),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1172 (.A(net1173),
    .X(net1172),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1173 (.A(_01516_),
    .X(net1173),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1174 (.A(_01435_),
    .X(net1174),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1175 (.A(net1179),
    .X(net1175),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1176 (.A(net1179),
    .X(net1176),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1177 (.A(net1178),
    .X(net1177),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1178 (.A(net1179),
    .X(net1178),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1179 (.A(\i_exotiny._0000_ ),
    .X(net1179),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1180 (.A(_01707_),
    .X(net1180),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1181 (.A(net1183),
    .X(net1181),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1182 (.A(net1183),
    .X(net1182),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1183 (.A(_01515_),
    .X(net1183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1184 (.A(_01472_),
    .X(net1184),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1185 (.A(net1187),
    .X(net1185),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1186 (.A(net1187),
    .X(net1186),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1187 (.A(_01451_),
    .X(net1187),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1188 (.A(net1189),
    .X(net1188),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1189 (.A(_01450_),
    .X(net1189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1190 (.A(net1191),
    .X(net1190),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1191 (.A(net1192),
    .X(net1191),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1192 (.A(net1193),
    .X(net1192),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1193 (.A(_01450_),
    .X(net1193),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1194 (.A(net1195),
    .X(net1194),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1195 (.A(net1197),
    .X(net1195),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1196 (.A(net1197),
    .X(net1196),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1197 (.A(net1200),
    .X(net1197),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1198 (.A(net1199),
    .X(net1198),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1199 (.A(net1200),
    .X(net1199),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1200 (.A(net3242),
    .X(net1200),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1201 (.A(_01434_),
    .X(net1201),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1202 (.A(_01434_),
    .X(net1202),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1203 (.A(\i_exotiny.i_wdg_top.cntr_inst.rst_n_sync ),
    .X(net1203),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1204 (.A(net1206),
    .X(net1204),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1205 (.A(net1206),
    .X(net1205),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1206 (.A(_02256_),
    .X(net1206),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1207 (.A(net1209),
    .X(net1207),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1208 (.A(net1209),
    .X(net1208),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1209 (.A(net1210),
    .X(net1209),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1210 (.A(net1211),
    .X(net1210),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1211 (.A(net1212),
    .X(net1211),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1212 (.A(_01504_),
    .X(net1212),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1213 (.A(net1217),
    .X(net1213),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1214 (.A(net1217),
    .X(net1214),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1215 (.A(net1217),
    .X(net1215),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1216 (.A(net1217),
    .X(net1216),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1217 (.A(_01503_),
    .X(net1217),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1218 (.A(_01489_),
    .X(net1218),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1219 (.A(_01447_),
    .X(net1219),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1220 (.A(net1221),
    .X(net1220),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1221 (.A(_01395_),
    .X(net1221),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1222 (.A(net1223),
    .X(net1222),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1223 (.A(_01394_),
    .X(net1223),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1224 (.A(_01382_),
    .X(net1224),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1225 (.A(net1226),
    .X(net1225),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1226 (.A(net1227),
    .X(net1226),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1227 (.A(_01378_),
    .X(net1227),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1228 (.A(net3839),
    .X(net1228),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1229 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[19] ),
    .X(net1229),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1230 (.A(net3699),
    .X(net1230),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1231 (.A(net1232),
    .X(net1231),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1232 (.A(net3732),
    .X(net1232),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1233 (.A(\i_exotiny._0315_[2] ),
    .X(net1233),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1234 (.A(net3688),
    .X(net1234),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1235 (.A(net1237),
    .X(net1235),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1236 (.A(net1237),
    .X(net1236),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1237 (.A(\i_exotiny._0079_[4] ),
    .X(net1237),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1238 (.A(net1239),
    .X(net1238),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1239 (.A(net3836),
    .X(net1239),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1240 (.A(net1241),
    .X(net1240),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1241 (.A(net3837),
    .X(net1241),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1242 (.A(\i_exotiny._0571_ ),
    .X(net1242),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1243 (.A(\i_exotiny._0601_ ),
    .X(net1243),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1244 (.A(net3767),
    .X(net1244),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1245 (.A(\i_exotiny._0542_ ),
    .X(net1245),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1246 (.A(net3807),
    .X(net1246),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1247 (.A(\i_exotiny._0590_ ),
    .X(net1247),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1248 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[5] ),
    .X(net1248),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1249 (.A(net3813),
    .X(net1249),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1250 (.A(net1251),
    .X(net1250),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1251 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[4] ),
    .X(net1251),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1252 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[3] ),
    .X(net1252),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1253 (.A(net1254),
    .X(net1253),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1254 (.A(net3469),
    .X(net1254),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1255 (.A(net1257),
    .X(net1255),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1256 (.A(net1257),
    .X(net1256),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1257 (.A(net3831),
    .X(net1257),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1258 (.A(net1259),
    .X(net1258),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1259 (.A(net3812),
    .X(net1259),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1260 (.A(net1261),
    .X(net1260),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1261 (.A(net3804),
    .X(net1261),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1262 (.A(net3144),
    .X(net1262),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1263 (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_hw_set [0]),
    .X(net1263),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1264 (.A(net3815),
    .X(net1264),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1265 (.A(net3833),
    .X(net1265),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1266 (.A(net1267),
    .X(net1266),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1267 (.A(net3694),
    .X(net1267),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1268 (.A(net3840),
    .X(net1268),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1269 (.A(net3840),
    .X(net1269),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1270 (.A(net3754),
    .X(net1270),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1271 (.A(net1274),
    .X(net1271),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1272 (.A(net1274),
    .X(net1272),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1273 (.A(net1274),
    .X(net1273),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1274 (.A(\i_exotiny._1312_ ),
    .X(net1274),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1275 (.A(net1278),
    .X(net1275),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1276 (.A(net1277),
    .X(net1276),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1277 (.A(net1278),
    .X(net1277),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1278 (.A(net1280),
    .X(net1278),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1279 (.A(net1280),
    .X(net1279),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1280 (.A(\i_exotiny._1312_ ),
    .X(net1280),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1281 (.A(net1282),
    .X(net1281),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1282 (.A(net1291),
    .X(net1282),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1283 (.A(net1285),
    .X(net1283),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1284 (.A(net1285),
    .X(net1284),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1285 (.A(net1291),
    .X(net1285),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1286 (.A(net1287),
    .X(net1286),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1287 (.A(net1289),
    .X(net1287),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout1288 (.A(net1289),
    .X(net1288),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1289 (.A(net1290),
    .X(net1289),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout1290 (.A(net1291),
    .X(net1290),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout1291 (.A(net3571),
    .X(net1291),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input10 (.A(uio_in[0]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input11 (.A(uio_in[1]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input12 (.A(uio_in[2]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input13 (.A(uio_in[3]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input14 (.A(uio_in[4]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(uio_in[5]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input16 (.A(uio_in[6]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input17 (.A(uio_in[7]),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_oe[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uio_oe[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uio_oe[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uio_oe[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uio_oe[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uio_oe[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uio_oe[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uio_oe[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uio_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output27 (.A(net27),
    .X(uio_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output28 (.A(net28),
    .X(uio_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output29 (.A(net29),
    .X(uio_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output30 (.A(net30),
    .X(uio_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output31 (.A(net31),
    .X(uio_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output32 (.A(net32),
    .X(uio_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output33 (.A(net33),
    .X(uio_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output34 (.A(net34),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output35 (.A(net35),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output36 (.A(net36),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output37 (.A(net37),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output38 (.A(net38),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output39 (.A(net39),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output40 (.A(net40),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output41 (.A(net41),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tiehi _09286__42 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net42));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_0_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_1_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_20_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_30_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_31_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_33_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_36_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_37_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_38_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_38_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_39_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_39_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_40_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_40_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_41_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_41_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_42_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_42_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_43_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_43_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_44_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_44_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_45_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_45_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_46_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_46_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_48_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_48_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_49_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_49_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_50_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_50_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_51_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_51_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_52_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_52_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_53_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_53_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_54_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_54_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_55_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_55_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_56_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_56_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_57_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_57_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_58_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_58_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_59_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_59_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_60_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_60_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_61_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_61_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_62_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_62_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_63_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_63_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_64_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_64_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_65_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_65_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_66_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_66_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_67_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_67_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_68_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_68_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_69_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_69_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_70_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_70_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_71_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_71_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_72_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_72_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_73_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_73_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_74_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_74_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_75_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_75_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_76_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_76_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_77_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_77_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_78_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_78_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_79_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_79_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_80_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_80_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_81_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_81_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_82_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_82_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_83_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_83_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_84_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_84_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_85_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_85_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_86_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_86_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_87_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_87_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_89_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_89_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_90_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_90_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_91_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_91_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_92_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_92_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_93_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_93_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_94_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_94_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_95_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_95_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_96_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_96_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_97_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_97_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_98_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_98_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_99_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_99_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_100_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_100_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_101_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_101_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_102_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_102_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_103_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_103_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_104_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_104_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_105_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_105_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_106_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_106_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_107_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_107_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_108_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_108_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_109_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_109_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_110_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_110_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_111_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_111_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_112_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_112_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_113_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_113_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_114_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_114_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_115_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_115_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_116_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_116_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_117_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_117_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_118_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_118_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_119_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_119_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_120_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_120_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_121_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_121_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_122_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_122_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_123_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_123_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_124_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_124_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_125_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_125_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_126_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_126_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_127_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_127_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_128_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_128_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_129_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_129_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_130_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_130_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_131_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_131_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_132_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_132_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_133_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_133_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_134_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_134_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_135_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_135_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_136_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_136_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_137_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_137_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_138_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_138_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_139_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_139_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_140_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_140_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_141_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_141_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_142_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_142_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_143_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_143_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_144_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_144_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_145_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_145_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_146_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_146_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_147_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_147_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_148_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_148_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_149_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_149_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_150_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_150_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_151_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_151_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_152_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_152_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_153_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_153_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_154_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_154_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_155_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_155_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_156_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_156_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_157_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_157_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_158_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_158_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_159_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_159_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_160_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_160_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_161_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_161_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_162_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_162_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_163_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_163_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_164_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_164_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_165_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_165_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_166_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_166_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_167_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_167_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_168_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_168_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_169_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_169_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_170_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_170_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_171_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_171_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_172_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_172_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_173_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_173_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_174_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_174_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_175_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_175_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_176_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_176_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_177_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_177_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_178_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_178_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_179_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_179_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_180_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_180_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_181_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_181_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_182_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_182_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_183_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_183_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_184_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_184_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_185_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_185_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_186_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_186_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_0__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_1__f_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_2__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_3__f_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_4__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_5__f_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_6__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_7__f_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_8__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_9__f_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_10__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_11__f_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_12__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_13__f_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_14__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_15__f_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_16__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_17__f_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_18__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_19__f_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_20__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_21__f_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_22__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_23__f_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_24__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_25__f_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_26__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_27__f_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_28__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_29__f_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_30__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_31__f_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload0 (.A(clknet_5_2__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload1 (.A(clknet_5_7__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload2 (.A(clknet_5_11__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload3 (.A(clknet_5_15__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload4 (.A(clknet_5_23__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload5 (.A(clknet_5_27__leaf_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload6 (.VDD(VPWR),
    .A(clknet_5_31__leaf_clk_regs),
    .VSS(VGND));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_186_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload8 (.VDD(VPWR),
    .A(clknet_leaf_180_clk_regs),
    .VSS(VGND));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_4_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload10 (.A(clknet_leaf_6_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload11 (.A(clknet_leaf_10_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload12 (.VDD(VPWR),
    .A(clknet_leaf_11_clk_regs),
    .VSS(VGND));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_12_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_17_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_162_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload16 (.A(clknet_leaf_115_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_159_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload18 (.A(clknet_leaf_161_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_9_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload20 (.VDD(VPWR),
    .A(clknet_leaf_32_clk_regs),
    .VSS(VGND));
 sg13g2_inv_4 clkload21 (.A(clknet_leaf_26_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_27_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload23 (.A(clknet_leaf_28_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload24 (.A(clknet_leaf_36_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload25 (.A(clknet_leaf_45_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload26 (.A(clknet_leaf_21_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload27 (.VDD(VPWR),
    .A(clknet_leaf_24_clk_regs),
    .VSS(VGND));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_50_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload29 (.VDD(VPWR),
    .A(clknet_leaf_58_clk_regs),
    .VSS(VGND));
 sg13g2_inv_2 clkload30 (.A(clknet_leaf_51_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_145_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload32 (.A(clknet_leaf_138_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload33 (.VDD(VPWR),
    .A(clknet_leaf_156_clk_regs),
    .VSS(VGND));
 sg13g2_inv_1 clkload34 (.VDD(VPWR),
    .A(clknet_leaf_130_clk_regs),
    .VSS(VGND));
 sg13g2_inv_2 clkload35 (.A(clknet_leaf_136_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload36 (.VDD(VPWR),
    .A(clknet_leaf_137_clk_regs),
    .VSS(VGND));
 sg13g2_inv_1 clkload37 (.VDD(VPWR),
    .A(clknet_leaf_104_clk_regs),
    .VSS(VGND));
 sg13g2_inv_1 clkload38 (.VDD(VPWR),
    .A(clknet_leaf_124_clk_regs),
    .VSS(VGND));
 sg13g2_inv_1 clkload39 (.VDD(VPWR),
    .A(clknet_leaf_67_clk_regs),
    .VSS(VGND));
 sg13g2_buf_8 clkload40 (.A(clknet_leaf_82_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload41 (.VDD(VPWR),
    .A(clknet_leaf_106_clk_regs),
    .VSS(VGND));
 sg13g2_buf_8 clkload42 (.A(clknet_leaf_89_clk_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload43 (.VDD(VPWR),
    .A(clknet_leaf_91_clk_regs),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1828));
 sg13g2_dlygate4sd3_1 hold2 (.A(_00804_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1829));
 sg13g2_dlygate4sd3_1 hold3 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1830));
 sg13g2_dlygate4sd3_1 hold4 (.A(_01115_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1831));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i_exotiny.i_wdg_top.fsm_inst.sw_trg_s1wto ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1832));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_exotiny._2055_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1833));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_exotiny.i_wb_spi.state_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1834));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_exotiny.i_wb_spi.state_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1835));
 sg13g2_dlygate4sd3_1 hold9 (.A(_00873_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1836));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_exotiny.i_wb_spi.state_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1837));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_exotiny.i_wb_spi.state_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1838));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_exotiny.i_wb_spi.state_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1839));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_exotiny.i_wb_spi.cnt_presc_r[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1840));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_exotiny.i_wb_spi.state_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1841));
 sg13g2_dlygate4sd3_1 hold15 (.A(_00874_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1842));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_exotiny.i_wb_spi.state_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1843));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_exotiny.i_wb_spi.state_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1844));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_exotiny.i_wb_spi.state_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1845));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_exotiny.i_wb_spi.state_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1846));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_exotiny.i_wb_spi.state_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1847));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_exotiny.i_wb_spi.state_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1848));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_exotiny.i_wb_spi.state_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1849));
 sg13g2_dlygate4sd3_1 hold23 (.A(_00871_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1850));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_exotiny.i_wb_spi.state_r[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1851));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_exotiny.i_wb_spi.state_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1852));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_exotiny.i_wb_spi.state_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1853));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i_exotiny.i_wb_spi.state_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1854));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_exotiny.i_wb_spi.state_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1855));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i_exotiny.i_wb_spi.state_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1856));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_exotiny.i_wb_spi.state_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1857));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_exotiny.i_wb_spi.state_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1858));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_exotiny.i_wb_spi.state_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1859));
 sg13g2_dlygate4sd3_1 hold33 (.A(_00876_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1860));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_exotiny.i_wb_spi.state_r[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1861));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_exotiny.i_wb_spi.state_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1862));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_exotiny.i_wb_spi.state_r[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1863));
 sg13g2_dlygate4sd3_1 hold37 (.A(\i_exotiny.i_wb_spi.state_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1864));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_exotiny.i_wb_spi.state_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1865));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_exotiny.i_wb_spi.state_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1866));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_exotiny.i_wb_spi.state_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1867));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_exotiny.i_wb_spi.state_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1868));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_exotiny.i_wb_spi.state_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1869));
 sg13g2_dlygate4sd3_1 hold43 (.A(\i_exotiny.i_wdg_top.o_wb_dat[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1870));
 sg13g2_dlygate4sd3_1 hold44 (.A(_00077_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1871));
 sg13g2_dlygate4sd3_1 hold45 (.A(\i_exotiny._0369_[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1872));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_exotiny.i_wdg_top.o_wb_dat[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1873));
 sg13g2_dlygate4sd3_1 hold47 (.A(_00079_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1874));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_exotiny.i_wdg_top.o_wb_dat[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1875));
 sg13g2_dlygate4sd3_1 hold49 (.A(_00078_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1876));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1877));
 sg13g2_dlygate4sd3_1 hold51 (.A(_03169_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1878));
 sg13g2_dlygate4sd3_1 hold52 (.A(_01125_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1879));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1880));
 sg13g2_dlygate4sd3_1 hold54 (.A(_03179_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1881));
 sg13g2_dlygate4sd3_1 hold55 (.A(_01131_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1882));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_exotiny.i_rstctl.cnt[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1883));
 sg13g2_dlygate4sd3_1 hold57 (.A(_01105_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1884));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1885));
 sg13g2_dlygate4sd3_1 hold59 (.A(_03157_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1886));
 sg13g2_dlygate4sd3_1 hold60 (.A(_01118_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1887));
 sg13g2_dlygate4sd3_1 hold61 (.A(_00020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1888));
 sg13g2_dlygate4sd3_1 hold62 (.A(_00076_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1889));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1890));
 sg13g2_dlygate4sd3_1 hold64 (.A(_03172_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1891));
 sg13g2_dlygate4sd3_1 hold65 (.A(_01127_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1892));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_exotiny._1429_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1893));
 sg13g2_dlygate4sd3_1 hold67 (.A(_01495_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1894));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_exotiny._1924_[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1895));
 sg13g2_dlygate4sd3_1 hold69 (.A(_00032_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1896));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_exotiny.i_wb_spi.dat_rx_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1897));
 sg13g2_dlygate4sd3_1 hold71 (.A(_00940_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1898));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_exotiny._1924_[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1899));
 sg13g2_dlygate4sd3_1 hold73 (.A(_00054_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1900));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_exotiny._1924_[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1901));
 sg13g2_dlygate4sd3_1 hold75 (.A(_00043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1902));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_exotiny._1924_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1903));
 sg13g2_dlygate4sd3_1 hold77 (.A(_00028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1904));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_exotiny.i_wb_spi.dat_rx_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1905));
 sg13g2_dlygate4sd3_1 hold79 (.A(_00941_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1906));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_exotiny._1924_[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1907));
 sg13g2_dlygate4sd3_1 hold81 (.A(_00029_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1908));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_exotiny._1924_[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1909));
 sg13g2_dlygate4sd3_1 hold83 (.A(_00036_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1910));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_exotiny._1160_[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1911));
 sg13g2_dlygate4sd3_1 hold85 (.A(_01064_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1912));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1913));
 sg13g2_dlygate4sd3_1 hold87 (.A(_03162_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1914));
 sg13g2_dlygate4sd3_1 hold88 (.A(_01121_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1915));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_exotiny._1924_[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1916));
 sg13g2_dlygate4sd3_1 hold90 (.A(_00046_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1917));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_exotiny._1924_[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1918));
 sg13g2_dlygate4sd3_1 hold92 (.A(_00053_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1919));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_exotiny._1924_[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1920));
 sg13g2_dlygate4sd3_1 hold94 (.A(_00050_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1921));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_exotiny._1924_[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1922));
 sg13g2_dlygate4sd3_1 hold96 (.A(_00037_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1923));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_exotiny._1924_[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1924));
 sg13g2_dlygate4sd3_1 hold98 (.A(_00052_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1925));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_exotiny._1924_[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1926));
 sg13g2_dlygate4sd3_1 hold100 (.A(_00047_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1927));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_exotiny.i_wb_spi.spi_sdo_o ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1928));
 sg13g2_dlygate4sd3_1 hold102 (.A(_00057_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1929));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1930));
 sg13g2_dlygate4sd3_1 hold104 (.A(_02380_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1931));
 sg13g2_dlygate4sd3_1 hold105 (.A(_00061_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1932));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_exotiny.i_wb_spi.dat_rx_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1933));
 sg13g2_dlygate4sd3_1 hold107 (.A(_00937_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1934));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_exotiny.i_wb_spi.dat_rx_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1935));
 sg13g2_dlygate4sd3_1 hold109 (.A(_00935_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1936));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_exotiny.i_wb_spi.dat_rx_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1937));
 sg13g2_dlygate4sd3_1 hold111 (.A(_00946_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1938));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_exotiny._1924_[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1939));
 sg13g2_dlygate4sd3_1 hold113 (.A(_00039_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1940));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_exotiny._1924_[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1941));
 sg13g2_dlygate4sd3_1 hold115 (.A(_00033_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1942));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_exotiny._1924_[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1943));
 sg13g2_dlygate4sd3_1 hold117 (.A(_00034_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1944));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_exotiny.i_wb_spi.dat_rx_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1945));
 sg13g2_dlygate4sd3_1 hold119 (.A(_00942_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1946));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_exotiny._1924_[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1947));
 sg13g2_dlygate4sd3_1 hold121 (.A(_00044_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1948));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_exotiny._1160_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1949));
 sg13g2_dlygate4sd3_1 hold123 (.A(_01040_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1950));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_exotiny.i_wb_spi.dat_rx_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1951));
 sg13g2_dlygate4sd3_1 hold125 (.A(_00945_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1952));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_exotiny._1924_[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1953));
 sg13g2_dlygate4sd3_1 hold127 (.A(_00038_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1954));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_exotiny._1160_[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1955));
 sg13g2_dlygate4sd3_1 hold129 (.A(_01044_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1956));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_exotiny._1924_[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1957));
 sg13g2_dlygate4sd3_1 hold131 (.A(_00045_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1958));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_exotiny._1924_[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1959));
 sg13g2_dlygate4sd3_1 hold133 (.A(_00056_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1960));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_exotiny._1924_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1961));
 sg13g2_dlygate4sd3_1 hold135 (.A(_01232_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1962));
 sg13g2_dlygate4sd3_1 hold136 (.A(\i_exotiny._1924_[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1963));
 sg13g2_dlygate4sd3_1 hold137 (.A(_00040_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1964));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_exotiny._0314_[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1965));
 sg13g2_dlygate4sd3_1 hold139 (.A(_00650_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1966));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_exotiny.i_wb_spi.dat_rx_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1967));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_exotiny.i_wb_spi.dat_rx_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1968));
 sg13g2_dlygate4sd3_1 hold142 (.A(_00936_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1969));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_exotiny.i_rstctl.cnt[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1970));
 sg13g2_dlygate4sd3_1 hold144 (.A(_01111_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1971));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1972));
 sg13g2_dlygate4sd3_1 hold146 (.A(_00059_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1973));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_exotiny._0314_[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1974));
 sg13g2_dlygate4sd3_1 hold148 (.A(_00651_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1975));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1976));
 sg13g2_dlygate4sd3_1 hold150 (.A(_00459_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1977));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_exotiny._1924_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1978));
 sg13g2_dlygate4sd3_1 hold152 (.A(_00027_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1979));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_exotiny._1612_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1980));
 sg13g2_dlygate4sd3_1 hold154 (.A(_00209_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1981));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_exotiny._1924_[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1982));
 sg13g2_dlygate4sd3_1 hold156 (.A(_00051_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1983));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1984));
 sg13g2_dlygate4sd3_1 hold158 (.A(_02254_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1985));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_exotiny._1489_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1986));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_exotiny._1924_[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1987));
 sg13g2_dlygate4sd3_1 hold161 (.A(_00031_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1988));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_exotiny._1160_[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1989));
 sg13g2_dlygate4sd3_1 hold163 (.A(_01041_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1990));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1991));
 sg13g2_dlygate4sd3_1 hold165 (.A(_02389_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1992));
 sg13g2_dlygate4sd3_1 hold166 (.A(_00065_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1993));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1994));
 sg13g2_dlygate4sd3_1 hold168 (.A(_00748_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1995));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_exotiny._1160_[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1996));
 sg13g2_dlygate4sd3_1 hold170 (.A(_01042_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1997));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_exotiny._1924_[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1998));
 sg13g2_dlygate4sd3_1 hold172 (.A(_00055_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1999));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2000));
 sg13g2_dlygate4sd3_1 hold174 (.A(_00462_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2001));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_exotiny._0314_[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2002));
 sg13g2_dlygate4sd3_1 hold176 (.A(_00657_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2003));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_exotiny._1924_[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2004));
 sg13g2_dlygate4sd3_1 hold178 (.A(_00041_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2005));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_exotiny._1924_[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2006));
 sg13g2_dlygate4sd3_1 hold180 (.A(_00035_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2007));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_exotiny._0314_[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2008));
 sg13g2_dlygate4sd3_1 hold182 (.A(_00649_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2009));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_exotiny._1160_[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2010));
 sg13g2_dlygate4sd3_1 hold184 (.A(_01050_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2011));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_exotiny._1614_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2012));
 sg13g2_dlygate4sd3_1 hold186 (.A(_00216_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2013));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_exotiny._0369_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2014));
 sg13g2_dlygate4sd3_1 hold188 (.A(_00514_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2015));
 sg13g2_dlygate4sd3_1 hold189 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2016));
 sg13g2_dlygate4sd3_1 hold190 (.A(_00465_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2017));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2018));
 sg13g2_dlygate4sd3_1 hold192 (.A(_00236_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2019));
 sg13g2_dlygate4sd3_1 hold193 (.A(\i_exotiny._1160_[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2020));
 sg13g2_dlygate4sd3_1 hold194 (.A(_01052_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2021));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_exotiny._1160_[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2022));
 sg13g2_dlygate4sd3_1 hold196 (.A(_01045_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2023));
 sg13g2_dlygate4sd3_1 hold197 (.A(\i_exotiny._0315_[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2024));
 sg13g2_dlygate4sd3_1 hold198 (.A(_01101_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2025));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_exotiny._1160_[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2026));
 sg13g2_dlygate4sd3_1 hold200 (.A(_01043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2027));
 sg13g2_dlygate4sd3_1 hold201 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2028));
 sg13g2_dlygate4sd3_1 hold202 (.A(_03164_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2029));
 sg13g2_dlygate4sd3_1 hold203 (.A(_01122_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2030));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_exotiny._1924_[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2031));
 sg13g2_dlygate4sd3_1 hold205 (.A(_00042_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2032));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.genblk7.g_value.r_value [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2033));
 sg13g2_dlygate4sd3_1 hold207 (.A(_00058_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2034));
 sg13g2_dlygate4sd3_1 hold208 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2035));
 sg13g2_dlygate4sd3_1 hold209 (.A(_01006_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2036));
 sg13g2_dlygate4sd3_1 hold210 (.A(\i_exotiny._0314_[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2037));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_exotiny._0314_[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2038));
 sg13g2_dlygate4sd3_1 hold212 (.A(_00648_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2039));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_exotiny._1160_[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2040));
 sg13g2_dlygate4sd3_1 hold214 (.A(_01051_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2041));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_exotiny._1615_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2042));
 sg13g2_dlygate4sd3_1 hold216 (.A(_00211_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2043));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_exotiny._1160_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2044));
 sg13g2_dlygate4sd3_1 hold218 (.A(_01038_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2045));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_exotiny._1924_[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2046));
 sg13g2_dlygate4sd3_1 hold220 (.A(_00048_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2047));
 sg13g2_dlygate4sd3_1 hold221 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2048));
 sg13g2_dlygate4sd3_1 hold222 (.A(_01219_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2049));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_exotiny._1924_[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2050));
 sg13g2_dlygate4sd3_1 hold224 (.A(_00030_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2051));
 sg13g2_dlygate4sd3_1 hold225 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2052));
 sg13g2_dlygate4sd3_1 hold226 (.A(_00909_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2053));
 sg13g2_dlygate4sd3_1 hold227 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2054));
 sg13g2_dlygate4sd3_1 hold228 (.A(_03181_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2055));
 sg13g2_dlygate4sd3_1 hold229 (.A(_01132_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2056));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2057));
 sg13g2_dlygate4sd3_1 hold231 (.A(_00529_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2058));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2059));
 sg13g2_dlygate4sd3_1 hold233 (.A(_00763_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2060));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_exotiny._0369_[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2061));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_exotiny._1611_[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2062));
 sg13g2_dlygate4sd3_1 hold236 (.A(\i_exotiny._1614_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2063));
 sg13g2_dlygate4sd3_1 hold237 (.A(_00215_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2064));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_exotiny._1160_[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2065));
 sg13g2_dlygate4sd3_1 hold239 (.A(_01046_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2066));
 sg13g2_dlygate4sd3_1 hold240 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2067));
 sg13g2_dlygate4sd3_1 hold241 (.A(_01001_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2068));
 sg13g2_dlygate4sd3_1 hold242 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2069));
 sg13g2_dlygate4sd3_1 hold243 (.A(_01329_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2070));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2071));
 sg13g2_dlygate4sd3_1 hold245 (.A(_01269_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2072));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2073));
 sg13g2_dlygate4sd3_1 hold247 (.A(_00265_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2074));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2075));
 sg13g2_dlygate4sd3_1 hold249 (.A(_00776_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2076));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_exotiny._1160_[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2077));
 sg13g2_dlygate4sd3_1 hold251 (.A(_01049_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2078));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2079));
 sg13g2_dlygate4sd3_1 hold253 (.A(_00894_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2080));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2081));
 sg13g2_dlygate4sd3_1 hold255 (.A(_00557_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2082));
 sg13g2_dlygate4sd3_1 hold256 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2083));
 sg13g2_dlygate4sd3_1 hold257 (.A(_00787_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2084));
 sg13g2_dlygate4sd3_1 hold258 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2085));
 sg13g2_dlygate4sd3_1 hold259 (.A(_00084_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2086));
 sg13g2_dlygate4sd3_1 hold260 (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.genblk7.g_value.r_value [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2087));
 sg13g2_dlygate4sd3_1 hold261 (.A(_00346_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2088));
 sg13g2_dlygate4sd3_1 hold262 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2089));
 sg13g2_dlygate4sd3_1 hold263 (.A(_00768_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2090));
 sg13g2_dlygate4sd3_1 hold264 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2091));
 sg13g2_dlygate4sd3_1 hold265 (.A(_00107_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2092));
 sg13g2_dlygate4sd3_1 hold266 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2093));
 sg13g2_dlygate4sd3_1 hold267 (.A(_00766_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2094));
 sg13g2_dlygate4sd3_1 hold268 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2095));
 sg13g2_dlygate4sd3_1 hold269 (.A(_00379_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2096));
 sg13g2_dlygate4sd3_1 hold270 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2097));
 sg13g2_dlygate4sd3_1 hold271 (.A(_01139_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2098));
 sg13g2_dlygate4sd3_1 hold272 (.A(\i_exotiny._0315_[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2099));
 sg13g2_dlygate4sd3_1 hold273 (.A(_01098_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2100));
 sg13g2_dlygate4sd3_1 hold274 (.A(\i_exotiny._1160_[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2101));
 sg13g2_dlygate4sd3_1 hold275 (.A(_01047_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2102));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2103));
 sg13g2_dlygate4sd3_1 hold277 (.A(_01013_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2104));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_exotiny.i_wb_spi.dat_rx_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2105));
 sg13g2_dlygate4sd3_1 hold279 (.A(\i_exotiny.i_wb_regs.spi_cpol_o ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2106));
 sg13g2_dlygate4sd3_1 hold280 (.A(_02955_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2107));
 sg13g2_dlygate4sd3_1 hold281 (.A(_00924_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2108));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2109));
 sg13g2_dlygate4sd3_1 hold283 (.A(_00330_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2110));
 sg13g2_dlygate4sd3_1 hold284 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2111));
 sg13g2_dlygate4sd3_1 hold285 (.A(_00785_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2112));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2113));
 sg13g2_dlygate4sd3_1 hold287 (.A(_00460_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2114));
 sg13g2_dlygate4sd3_1 hold288 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2115));
 sg13g2_dlygate4sd3_1 hold289 (.A(_00285_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2116));
 sg13g2_dlygate4sd3_1 hold290 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2117));
 sg13g2_dlygate4sd3_1 hold291 (.A(_00846_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2118));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2119));
 sg13g2_dlygate4sd3_1 hold293 (.A(_00412_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2120));
 sg13g2_dlygate4sd3_1 hold294 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2121));
 sg13g2_dlygate4sd3_1 hold295 (.A(_01323_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2122));
 sg13g2_dlygate4sd3_1 hold296 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2123));
 sg13g2_dlygate4sd3_1 hold297 (.A(_00130_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2124));
 sg13g2_dlygate4sd3_1 hold298 (.A(\i_exotiny._0369_[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2125));
 sg13g2_dlygate4sd3_1 hold299 (.A(\i_exotiny._1611_[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2126));
 sg13g2_dlygate4sd3_1 hold300 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2127));
 sg13g2_dlygate4sd3_1 hold301 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2128));
 sg13g2_dlygate4sd3_1 hold302 (.A(_00113_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2129));
 sg13g2_dlygate4sd3_1 hold303 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2130));
 sg13g2_dlygate4sd3_1 hold304 (.A(_01153_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2131));
 sg13g2_dlygate4sd3_1 hold305 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2132));
 sg13g2_dlygate4sd3_1 hold306 (.A(_01255_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2133));
 sg13g2_dlygate4sd3_1 hold307 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2134));
 sg13g2_dlygate4sd3_1 hold308 (.A(_01297_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2135));
 sg13g2_dlygate4sd3_1 hold309 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2136));
 sg13g2_dlygate4sd3_1 hold310 (.A(_00382_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2137));
 sg13g2_dlygate4sd3_1 hold311 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2138));
 sg13g2_dlygate4sd3_1 hold312 (.A(_00475_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2139));
 sg13g2_dlygate4sd3_1 hold313 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2140));
 sg13g2_dlygate4sd3_1 hold314 (.A(_00249_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2141));
 sg13g2_dlygate4sd3_1 hold315 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2142));
 sg13g2_dlygate4sd3_1 hold316 (.A(_01307_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2143));
 sg13g2_dlygate4sd3_1 hold317 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2144));
 sg13g2_dlygate4sd3_1 hold318 (.A(_00836_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2145));
 sg13g2_dlygate4sd3_1 hold319 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2146));
 sg13g2_dlygate4sd3_1 hold320 (.A(_00347_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2147));
 sg13g2_dlygate4sd3_1 hold321 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2148));
 sg13g2_dlygate4sd3_1 hold322 (.A(_00259_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2149));
 sg13g2_dlygate4sd3_1 hold323 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2150));
 sg13g2_dlygate4sd3_1 hold324 (.A(_00611_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2151));
 sg13g2_dlygate4sd3_1 hold325 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2152));
 sg13g2_dlygate4sd3_1 hold326 (.A(_00092_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2153));
 sg13g2_dlygate4sd3_1 hold327 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2154));
 sg13g2_dlygate4sd3_1 hold328 (.A(_00184_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2155));
 sg13g2_dlygate4sd3_1 hold329 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2156));
 sg13g2_dlygate4sd3_1 hold330 (.A(_00202_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2157));
 sg13g2_dlygate4sd3_1 hold331 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2158));
 sg13g2_dlygate4sd3_1 hold332 (.A(_00844_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2159));
 sg13g2_dlygate4sd3_1 hold333 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2160));
 sg13g2_dlygate4sd3_1 hold334 (.A(_00757_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2161));
 sg13g2_dlygate4sd3_1 hold335 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2162));
 sg13g2_dlygate4sd3_1 hold336 (.A(_01299_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2163));
 sg13g2_dlygate4sd3_1 hold337 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2164));
 sg13g2_dlygate4sd3_1 hold338 (.A(_00133_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2165));
 sg13g2_dlygate4sd3_1 hold339 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2166));
 sg13g2_dlygate4sd3_1 hold340 (.A(_00316_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2167));
 sg13g2_dlygate4sd3_1 hold341 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2168));
 sg13g2_dlygate4sd3_1 hold342 (.A(_00146_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2169));
 sg13g2_dlygate4sd3_1 hold343 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2170));
 sg13g2_dlygate4sd3_1 hold344 (.A(_00157_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2171));
 sg13g2_dlygate4sd3_1 hold345 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2172));
 sg13g2_dlygate4sd3_1 hold346 (.A(_01193_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2173));
 sg13g2_dlygate4sd3_1 hold347 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2174));
 sg13g2_dlygate4sd3_1 hold348 (.A(_00891_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2175));
 sg13g2_dlygate4sd3_1 hold349 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2176));
 sg13g2_dlygate4sd3_1 hold350 (.A(_01186_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2177));
 sg13g2_dlygate4sd3_1 hold351 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2178));
 sg13g2_dlygate4sd3_1 hold352 (.A(_00758_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2179));
 sg13g2_dlygate4sd3_1 hold353 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2180));
 sg13g2_dlygate4sd3_1 hold354 (.A(_00397_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2181));
 sg13g2_dlygate4sd3_1 hold355 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2182));
 sg13g2_dlygate4sd3_1 hold356 (.A(_01167_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2183));
 sg13g2_dlygate4sd3_1 hold357 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2184));
 sg13g2_dlygate4sd3_1 hold358 (.A(_00600_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2185));
 sg13g2_dlygate4sd3_1 hold359 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2186));
 sg13g2_dlygate4sd3_1 hold360 (.A(_01136_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2187));
 sg13g2_dlygate4sd3_1 hold361 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2188));
 sg13g2_dlygate4sd3_1 hold362 (.A(_01340_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2189));
 sg13g2_dlygate4sd3_1 hold363 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2190));
 sg13g2_dlygate4sd3_1 hold364 (.A(_01352_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2191));
 sg13g2_dlygate4sd3_1 hold365 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2192));
 sg13g2_dlygate4sd3_1 hold366 (.A(_00719_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2193));
 sg13g2_dlygate4sd3_1 hold367 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2194));
 sg13g2_dlygate4sd3_1 hold368 (.A(_01184_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2195));
 sg13g2_dlygate4sd3_1 hold369 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2196));
 sg13g2_dlygate4sd3_1 hold370 (.A(_00497_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2197));
 sg13g2_dlygate4sd3_1 hold371 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2198));
 sg13g2_dlygate4sd3_1 hold372 (.A(_00904_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2199));
 sg13g2_dlygate4sd3_1 hold373 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2200));
 sg13g2_dlygate4sd3_1 hold374 (.A(_00399_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2201));
 sg13g2_dlygate4sd3_1 hold375 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2202));
 sg13g2_dlygate4sd3_1 hold376 (.A(_00995_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2203));
 sg13g2_dlygate4sd3_1 hold377 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2204));
 sg13g2_dlygate4sd3_1 hold378 (.A(_00892_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2205));
 sg13g2_dlygate4sd3_1 hold379 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2206));
 sg13g2_dlygate4sd3_1 hold380 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2207));
 sg13g2_dlygate4sd3_1 hold381 (.A(_00178_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2208));
 sg13g2_dlygate4sd3_1 hold382 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2209));
 sg13g2_dlygate4sd3_1 hold383 (.A(_01194_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2210));
 sg13g2_dlygate4sd3_1 hold384 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2211));
 sg13g2_dlygate4sd3_1 hold385 (.A(_01342_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2212));
 sg13g2_dlygate4sd3_1 hold386 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2213));
 sg13g2_dlygate4sd3_1 hold387 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2214));
 sg13g2_dlygate4sd3_1 hold388 (.A(_00083_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2215));
 sg13g2_dlygate4sd3_1 hold389 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2216));
 sg13g2_dlygate4sd3_1 hold390 (.A(_00854_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2217));
 sg13g2_dlygate4sd3_1 hold391 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2218));
 sg13g2_dlygate4sd3_1 hold392 (.A(_00323_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2219));
 sg13g2_dlygate4sd3_1 hold393 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2220));
 sg13g2_dlygate4sd3_1 hold394 (.A(_00233_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2221));
 sg13g2_dlygate4sd3_1 hold395 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2222));
 sg13g2_dlygate4sd3_1 hold396 (.A(_00812_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2223));
 sg13g2_dlygate4sd3_1 hold397 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2224));
 sg13g2_dlygate4sd3_1 hold398 (.A(_00601_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2225));
 sg13g2_dlygate4sd3_1 hold399 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2226));
 sg13g2_dlygate4sd3_1 hold400 (.A(_00335_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2227));
 sg13g2_dlygate4sd3_1 hold401 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2228));
 sg13g2_dlygate4sd3_1 hold402 (.A(_00574_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2229));
 sg13g2_dlygate4sd3_1 hold403 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2230));
 sg13g2_dlygate4sd3_1 hold404 (.A(_00348_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2231));
 sg13g2_dlygate4sd3_1 hold405 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2232));
 sg13g2_dlygate4sd3_1 hold406 (.A(_00531_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2233));
 sg13g2_dlygate4sd3_1 hold407 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2234));
 sg13g2_dlygate4sd3_1 hold408 (.A(_00164_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2235));
 sg13g2_dlygate4sd3_1 hold409 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2236));
 sg13g2_dlygate4sd3_1 hold410 (.A(_01155_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2237));
 sg13g2_dlygate4sd3_1 hold411 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2238));
 sg13g2_dlygate4sd3_1 hold412 (.A(_00333_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2239));
 sg13g2_dlygate4sd3_1 hold413 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2240));
 sg13g2_dlygate4sd3_1 hold414 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2241));
 sg13g2_dlygate4sd3_1 hold415 (.A(_01246_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2242));
 sg13g2_dlygate4sd3_1 hold416 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2243));
 sg13g2_dlygate4sd3_1 hold417 (.A(_00733_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2244));
 sg13g2_dlygate4sd3_1 hold418 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2245));
 sg13g2_dlygate4sd3_1 hold419 (.A(_01008_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2246));
 sg13g2_dlygate4sd3_1 hold420 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2247));
 sg13g2_dlygate4sd3_1 hold421 (.A(_00094_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2248));
 sg13g2_dlygate4sd3_1 hold422 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2249));
 sg13g2_dlygate4sd3_1 hold423 (.A(_00547_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2250));
 sg13g2_dlygate4sd3_1 hold424 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2251));
 sg13g2_dlygate4sd3_1 hold425 (.A(_01276_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2252));
 sg13g2_dlygate4sd3_1 hold426 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2253));
 sg13g2_dlygate4sd3_1 hold427 (.A(_01353_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2254));
 sg13g2_dlygate4sd3_1 hold428 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2255));
 sg13g2_dlygate4sd3_1 hold429 (.A(_00252_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2256));
 sg13g2_dlygate4sd3_1 hold430 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2257));
 sg13g2_dlygate4sd3_1 hold431 (.A(_00237_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2258));
 sg13g2_dlygate4sd3_1 hold432 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2259));
 sg13g2_dlygate4sd3_1 hold433 (.A(_01347_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2260));
 sg13g2_dlygate4sd3_1 hold434 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2261));
 sg13g2_dlygate4sd3_1 hold435 (.A(_00300_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2262));
 sg13g2_dlygate4sd3_1 hold436 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2263));
 sg13g2_dlygate4sd3_1 hold437 (.A(_00329_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2264));
 sg13g2_dlygate4sd3_1 hold438 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2265));
 sg13g2_dlygate4sd3_1 hold439 (.A(_00712_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2266));
 sg13g2_dlygate4sd3_1 hold440 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2267));
 sg13g2_dlygate4sd3_1 hold441 (.A(_01324_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2268));
 sg13g2_dlygate4sd3_1 hold442 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2269));
 sg13g2_dlygate4sd3_1 hold443 (.A(_00482_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2270));
 sg13g2_dlygate4sd3_1 hold444 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2271));
 sg13g2_dlygate4sd3_1 hold445 (.A(_00243_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2272));
 sg13g2_dlygate4sd3_1 hold446 (.A(\i_exotiny._0022_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2273));
 sg13g2_dlygate4sd3_1 hold447 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2274));
 sg13g2_dlygate4sd3_1 hold448 (.A(_00589_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2275));
 sg13g2_dlygate4sd3_1 hold449 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2276));
 sg13g2_dlygate4sd3_1 hold450 (.A(_00274_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2277));
 sg13g2_dlygate4sd3_1 hold451 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2278));
 sg13g2_dlygate4sd3_1 hold452 (.A(_00717_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2279));
 sg13g2_dlygate4sd3_1 hold453 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2280));
 sg13g2_dlygate4sd3_1 hold454 (.A(_00746_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2281));
 sg13g2_dlygate4sd3_1 hold455 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2282));
 sg13g2_dlygate4sd3_1 hold456 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2283));
 sg13g2_dlygate4sd3_1 hold457 (.A(_00485_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2284));
 sg13g2_dlygate4sd3_1 hold458 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2285));
 sg13g2_dlygate4sd3_1 hold459 (.A(_00587_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2286));
 sg13g2_dlygate4sd3_1 hold460 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2287));
 sg13g2_dlygate4sd3_1 hold461 (.A(_00099_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2288));
 sg13g2_dlygate4sd3_1 hold462 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2289));
 sg13g2_dlygate4sd3_1 hold463 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2290));
 sg13g2_dlygate4sd3_1 hold464 (.A(_01018_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2291));
 sg13g2_dlygate4sd3_1 hold465 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2292));
 sg13g2_dlygate4sd3_1 hold466 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2293));
 sg13g2_dlygate4sd3_1 hold467 (.A(_00800_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2294));
 sg13g2_dlygate4sd3_1 hold468 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2295));
 sg13g2_dlygate4sd3_1 hold469 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2296));
 sg13g2_dlygate4sd3_1 hold470 (.A(_01165_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2297));
 sg13g2_dlygate4sd3_1 hold471 (.A(\i_exotiny.i_rstctl.cnt[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2298));
 sg13g2_dlygate4sd3_1 hold472 (.A(_03136_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2299));
 sg13g2_dlygate4sd3_1 hold473 (.A(_01107_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2300));
 sg13g2_dlygate4sd3_1 hold474 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2301));
 sg13g2_dlygate4sd3_1 hold475 (.A(_01176_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2302));
 sg13g2_dlygate4sd3_1 hold476 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2303));
 sg13g2_dlygate4sd3_1 hold477 (.A(_00253_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2304));
 sg13g2_dlygate4sd3_1 hold478 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2305));
 sg13g2_dlygate4sd3_1 hold479 (.A(_00372_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2306));
 sg13g2_dlygate4sd3_1 hold480 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2307));
 sg13g2_dlygate4sd3_1 hold481 (.A(_01300_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2308));
 sg13g2_dlygate4sd3_1 hold482 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2309));
 sg13g2_dlygate4sd3_1 hold483 (.A(_00976_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2310));
 sg13g2_dlygate4sd3_1 hold484 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2311));
 sg13g2_dlygate4sd3_1 hold485 (.A(_00972_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2312));
 sg13g2_dlygate4sd3_1 hold486 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2313));
 sg13g2_dlygate4sd3_1 hold487 (.A(_00821_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2314));
 sg13g2_dlygate4sd3_1 hold488 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2315));
 sg13g2_dlygate4sd3_1 hold489 (.A(_00718_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2316));
 sg13g2_dlygate4sd3_1 hold490 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2317));
 sg13g2_dlygate4sd3_1 hold491 (.A(_00283_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2318));
 sg13g2_dlygate4sd3_1 hold492 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2319));
 sg13g2_dlygate4sd3_1 hold493 (.A(_00148_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2320));
 sg13g2_dlygate4sd3_1 hold494 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2321));
 sg13g2_dlygate4sd3_1 hold495 (.A(_00085_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2322));
 sg13g2_dlygate4sd3_1 hold496 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2323));
 sg13g2_dlygate4sd3_1 hold497 (.A(_00903_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2324));
 sg13g2_dlygate4sd3_1 hold498 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2325));
 sg13g2_dlygate4sd3_1 hold499 (.A(_00455_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2326));
 sg13g2_dlygate4sd3_1 hold500 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2327));
 sg13g2_dlygate4sd3_1 hold501 (.A(_01345_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2328));
 sg13g2_dlygate4sd3_1 hold502 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2329));
 sg13g2_dlygate4sd3_1 hold503 (.A(_00745_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2330));
 sg13g2_dlygate4sd3_1 hold504 (.A(\i_exotiny._1612_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2331));
 sg13g2_dlygate4sd3_1 hold505 (.A(_00210_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2332));
 sg13g2_dlygate4sd3_1 hold506 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2333));
 sg13g2_dlygate4sd3_1 hold507 (.A(_00305_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2334));
 sg13g2_dlygate4sd3_1 hold508 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2335));
 sg13g2_dlygate4sd3_1 hold509 (.A(_01207_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2336));
 sg13g2_dlygate4sd3_1 hold510 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2337));
 sg13g2_dlygate4sd3_1 hold511 (.A(_00199_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2338));
 sg13g2_dlygate4sd3_1 hold512 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2339));
 sg13g2_dlygate4sd3_1 hold513 (.A(_00974_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2340));
 sg13g2_dlygate4sd3_1 hold514 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2341));
 sg13g2_dlygate4sd3_1 hold515 (.A(_00584_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2342));
 sg13g2_dlygate4sd3_1 hold516 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2343));
 sg13g2_dlygate4sd3_1 hold517 (.A(_00192_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2344));
 sg13g2_dlygate4sd3_1 hold518 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2345));
 sg13g2_dlygate4sd3_1 hold519 (.A(_01284_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2346));
 sg13g2_dlygate4sd3_1 hold520 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2347));
 sg13g2_dlygate4sd3_1 hold521 (.A(_01318_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2348));
 sg13g2_dlygate4sd3_1 hold522 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2349));
 sg13g2_dlygate4sd3_1 hold523 (.A(_01158_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2350));
 sg13g2_dlygate4sd3_1 hold524 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2351));
 sg13g2_dlygate4sd3_1 hold525 (.A(_00126_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2352));
 sg13g2_dlygate4sd3_1 hold526 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2353));
 sg13g2_dlygate4sd3_1 hold527 (.A(_00473_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2354));
 sg13g2_dlygate4sd3_1 hold528 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2355));
 sg13g2_dlygate4sd3_1 hold529 (.A(_00755_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2356));
 sg13g2_dlygate4sd3_1 hold530 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2357));
 sg13g2_dlygate4sd3_1 hold531 (.A(_00128_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2358));
 sg13g2_dlygate4sd3_1 hold532 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2359));
 sg13g2_dlygate4sd3_1 hold533 (.A(_00830_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2360));
 sg13g2_dlygate4sd3_1 hold534 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2361));
 sg13g2_dlygate4sd3_1 hold535 (.A(_00966_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2362));
 sg13g2_dlygate4sd3_1 hold536 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2363));
 sg13g2_dlygate4sd3_1 hold537 (.A(_00581_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2364));
 sg13g2_dlygate4sd3_1 hold538 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2365));
 sg13g2_dlygate4sd3_1 hold539 (.A(_01334_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2366));
 sg13g2_dlygate4sd3_1 hold540 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2367));
 sg13g2_dlygate4sd3_1 hold541 (.A(_00432_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2368));
 sg13g2_dlygate4sd3_1 hold542 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2369));
 sg13g2_dlygate4sd3_1 hold543 (.A(_00368_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2370));
 sg13g2_dlygate4sd3_1 hold544 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2371));
 sg13g2_dlygate4sd3_1 hold545 (.A(_01330_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2372));
 sg13g2_dlygate4sd3_1 hold546 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2373));
 sg13g2_dlygate4sd3_1 hold547 (.A(_00400_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2374));
 sg13g2_dlygate4sd3_1 hold548 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2375));
 sg13g2_dlygate4sd3_1 hold549 (.A(_00367_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2376));
 sg13g2_dlygate4sd3_1 hold550 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2377));
 sg13g2_dlygate4sd3_1 hold551 (.A(_00186_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2378));
 sg13g2_dlygate4sd3_1 hold552 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2379));
 sg13g2_dlygate4sd3_1 hold553 (.A(_01224_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2380));
 sg13g2_dlygate4sd3_1 hold554 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2381));
 sg13g2_dlygate4sd3_1 hold555 (.A(_00535_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2382));
 sg13g2_dlygate4sd3_1 hold556 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2383));
 sg13g2_dlygate4sd3_1 hold557 (.A(_00439_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2384));
 sg13g2_dlygate4sd3_1 hold558 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2385));
 sg13g2_dlygate4sd3_1 hold559 (.A(_00422_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2386));
 sg13g2_dlygate4sd3_1 hold560 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2387));
 sg13g2_dlygate4sd3_1 hold561 (.A(_01222_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2388));
 sg13g2_dlygate4sd3_1 hold562 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2389));
 sg13g2_dlygate4sd3_1 hold563 (.A(_00307_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2390));
 sg13g2_dlygate4sd3_1 hold564 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2391));
 sg13g2_dlygate4sd3_1 hold565 (.A(_00238_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2392));
 sg13g2_dlygate4sd3_1 hold566 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2393));
 sg13g2_dlygate4sd3_1 hold567 (.A(_00807_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2394));
 sg13g2_dlygate4sd3_1 hold568 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2395));
 sg13g2_dlygate4sd3_1 hold569 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2396));
 sg13g2_dlygate4sd3_1 hold570 (.A(_01156_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2397));
 sg13g2_dlygate4sd3_1 hold571 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2398));
 sg13g2_dlygate4sd3_1 hold572 (.A(_00989_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2399));
 sg13g2_dlygate4sd3_1 hold573 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2400));
 sg13g2_dlygate4sd3_1 hold574 (.A(_00275_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2401));
 sg13g2_dlygate4sd3_1 hold575 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2402));
 sg13g2_dlygate4sd3_1 hold576 (.A(_00415_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2403));
 sg13g2_dlygate4sd3_1 hold577 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2404));
 sg13g2_dlygate4sd3_1 hold578 (.A(_01241_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2405));
 sg13g2_dlygate4sd3_1 hold579 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2406));
 sg13g2_dlygate4sd3_1 hold580 (.A(_00162_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2407));
 sg13g2_dlygate4sd3_1 hold581 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2408));
 sg13g2_dlygate4sd3_1 hold582 (.A(_00701_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2409));
 sg13g2_dlygate4sd3_1 hold583 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2410));
 sg13g2_dlygate4sd3_1 hold584 (.A(_00795_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2411));
 sg13g2_dlygate4sd3_1 hold585 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2412));
 sg13g2_dlygate4sd3_1 hold586 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2413));
 sg13g2_dlygate4sd3_1 hold587 (.A(_00268_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2414));
 sg13g2_dlygate4sd3_1 hold588 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2415));
 sg13g2_dlygate4sd3_1 hold589 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2416));
 sg13g2_dlygate4sd3_1 hold590 (.A(_00384_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2417));
 sg13g2_dlygate4sd3_1 hold591 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2418));
 sg13g2_dlygate4sd3_1 hold592 (.A(_00149_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2419));
 sg13g2_dlygate4sd3_1 hold593 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2420));
 sg13g2_dlygate4sd3_1 hold594 (.A(_01179_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2421));
 sg13g2_dlygate4sd3_1 hold595 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2422));
 sg13g2_dlygate4sd3_1 hold596 (.A(_01213_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2423));
 sg13g2_dlygate4sd3_1 hold597 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2424));
 sg13g2_dlygate4sd3_1 hold598 (.A(_00440_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2425));
 sg13g2_dlygate4sd3_1 hold599 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2426));
 sg13g2_dlygate4sd3_1 hold600 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2427));
 sg13g2_dlygate4sd3_1 hold601 (.A(_00357_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2428));
 sg13g2_dlygate4sd3_1 hold602 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2429));
 sg13g2_dlygate4sd3_1 hold603 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2430));
 sg13g2_dlygate4sd3_1 hold604 (.A(_00143_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2431));
 sg13g2_dlygate4sd3_1 hold605 (.A(\i_exotiny.i_wb_spi.dat_rx_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2432));
 sg13g2_dlygate4sd3_1 hold606 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2433));
 sg13g2_dlygate4sd3_1 hold607 (.A(_00131_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2434));
 sg13g2_dlygate4sd3_1 hold608 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2435));
 sg13g2_dlygate4sd3_1 hold609 (.A(_00273_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2436));
 sg13g2_dlygate4sd3_1 hold610 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2437));
 sg13g2_dlygate4sd3_1 hold611 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2438));
 sg13g2_dlygate4sd3_1 hold612 (.A(_00992_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2439));
 sg13g2_dlygate4sd3_1 hold613 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2440));
 sg13g2_dlygate4sd3_1 hold614 (.A(_00183_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2441));
 sg13g2_dlygate4sd3_1 hold615 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2442));
 sg13g2_dlygate4sd3_1 hold616 (.A(_00914_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2443));
 sg13g2_dlygate4sd3_1 hold617 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2444));
 sg13g2_dlygate4sd3_1 hold618 (.A(_00141_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2445));
 sg13g2_dlygate4sd3_1 hold619 (.A(\i_exotiny._0314_[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2446));
 sg13g2_dlygate4sd3_1 hold620 (.A(_00656_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2447));
 sg13g2_dlygate4sd3_1 hold621 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2448));
 sg13g2_dlygate4sd3_1 hold622 (.A(_00570_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2449));
 sg13g2_dlygate4sd3_1 hold623 (.A(\i_exotiny._0034_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2450));
 sg13g2_dlygate4sd3_1 hold624 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2451));
 sg13g2_dlygate4sd3_1 hold625 (.A(_01331_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2452));
 sg13g2_dlygate4sd3_1 hold626 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2453));
 sg13g2_dlygate4sd3_1 hold627 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2454));
 sg13g2_dlygate4sd3_1 hold628 (.A(_00979_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2455));
 sg13g2_dlygate4sd3_1 hold629 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2456));
 sg13g2_dlygate4sd3_1 hold630 (.A(_00167_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2457));
 sg13g2_dlygate4sd3_1 hold631 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2458));
 sg13g2_dlygate4sd3_1 hold632 (.A(_00165_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2459));
 sg13g2_dlygate4sd3_1 hold633 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2460));
 sg13g2_dlygate4sd3_1 hold634 (.A(_01240_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2461));
 sg13g2_dlygate4sd3_1 hold635 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2462));
 sg13g2_dlygate4sd3_1 hold636 (.A(_01137_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2463));
 sg13g2_dlygate4sd3_1 hold637 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2464));
 sg13g2_dlygate4sd3_1 hold638 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2465));
 sg13g2_dlygate4sd3_1 hold639 (.A(_00444_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2466));
 sg13g2_dlygate4sd3_1 hold640 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2467));
 sg13g2_dlygate4sd3_1 hold641 (.A(_00967_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2468));
 sg13g2_dlygate4sd3_1 hold642 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2469));
 sg13g2_dlygate4sd3_1 hold643 (.A(_01317_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2470));
 sg13g2_dlygate4sd3_1 hold644 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2471));
 sg13g2_dlygate4sd3_1 hold645 (.A(_01325_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2472));
 sg13g2_dlygate4sd3_1 hold646 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2473));
 sg13g2_dlygate4sd3_1 hold647 (.A(_00496_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2474));
 sg13g2_dlygate4sd3_1 hold648 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2475));
 sg13g2_dlygate4sd3_1 hold649 (.A(_00366_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2476));
 sg13g2_dlygate4sd3_1 hold650 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2477));
 sg13g2_dlygate4sd3_1 hold651 (.A(_00174_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2478));
 sg13g2_dlygate4sd3_1 hold652 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2479));
 sg13g2_dlygate4sd3_1 hold653 (.A(_00371_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2480));
 sg13g2_dlygate4sd3_1 hold654 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2481));
 sg13g2_dlygate4sd3_1 hold655 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2482));
 sg13g2_dlygate4sd3_1 hold656 (.A(_00112_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2483));
 sg13g2_dlygate4sd3_1 hold657 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2484));
 sg13g2_dlygate4sd3_1 hold658 (.A(_00080_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2485));
 sg13g2_dlygate4sd3_1 hold659 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2486));
 sg13g2_dlygate4sd3_1 hold660 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2487));
 sg13g2_dlygate4sd3_1 hold661 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2488));
 sg13g2_dlygate4sd3_1 hold662 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2489));
 sg13g2_dlygate4sd3_1 hold663 (.A(_00129_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2490));
 sg13g2_dlygate4sd3_1 hold664 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2491));
 sg13g2_dlygate4sd3_1 hold665 (.A(_00617_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2492));
 sg13g2_dlygate4sd3_1 hold666 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2493));
 sg13g2_dlygate4sd3_1 hold667 (.A(_00491_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2494));
 sg13g2_dlygate4sd3_1 hold668 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2495));
 sg13g2_dlygate4sd3_1 hold669 (.A(_01019_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold670 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold671 (.A(_01292_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold672 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2499));
 sg13g2_dlygate4sd3_1 hold673 (.A(_01189_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2500));
 sg13g2_dlygate4sd3_1 hold674 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2501));
 sg13g2_dlygate4sd3_1 hold675 (.A(_00095_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2502));
 sg13g2_dlygate4sd3_1 hold676 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2503));
 sg13g2_dlygate4sd3_1 hold677 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2504));
 sg13g2_dlygate4sd3_1 hold678 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2505));
 sg13g2_dlygate4sd3_1 hold679 (.A(_00175_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2506));
 sg13g2_dlygate4sd3_1 hold680 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold681 (.A(_00423_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold682 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold683 (.A(_00142_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold684 (.A(\i_exotiny._0030_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold685 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold686 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold687 (.A(_00220_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold688 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold689 (.A(_00498_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold690 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold691 (.A(_01225_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold692 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold693 (.A(_01256_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold694 (.A(\i_exotiny._0025_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold695 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold696 (.A(_00506_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold697 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold698 (.A(_00700_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold699 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold700 (.A(_01187_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold701 (.A(\i_exotiny._1924_[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold702 (.A(_00049_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold703 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold704 (.A(_00560_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold705 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold706 (.A(_00583_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold707 (.A(\i_exotiny._0021_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold708 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold709 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold710 (.A(_01320_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold711 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold712 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold713 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold714 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold715 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold716 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold717 (.A(_00101_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold718 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold719 (.A(_01208_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold720 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold721 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold722 (.A(_00803_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold723 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold724 (.A(_00532_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold725 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold726 (.A(_00121_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold727 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold728 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold729 (.A(_00818_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold730 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold731 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold732 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold733 (.A(_01260_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold734 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold735 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold736 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold737 (.A(_00231_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold738 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold739 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold740 (.A(_00365_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold741 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold742 (.A(_01214_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold743 (.A(\i_exotiny.i_rstctl.wdg_res_n ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold744 (.A(_02914_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold745 (.A(_00698_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold746 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold747 (.A(_00816_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold748 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold749 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold750 (.A(_00504_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold751 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold752 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold753 (.A(_01212_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold754 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold755 (.A(_01247_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold756 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold757 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold758 (.A(_00998_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold759 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold760 (.A(_00181_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold761 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold762 (.A(_00245_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold763 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold764 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold765 (.A(\i_exotiny._0022_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold766 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold767 (.A(_00271_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold768 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold769 (.A(_00189_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold770 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold771 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold772 (.A(_00090_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold773 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold774 (.A(_01234_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold775 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold776 (.A(_00293_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold777 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold778 (.A(_00226_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold779 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold780 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold781 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold782 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold783 (.A(_00530_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold784 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold785 (.A(_00228_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold786 (.A(\i_exotiny._0027_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold787 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold788 (.A(_00990_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold789 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold790 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold791 (.A(_00610_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold792 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold793 (.A(_00264_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold794 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold795 (.A(_00395_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold796 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold797 (.A(_00607_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold798 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold799 (.A(_01282_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold800 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold801 (.A(_00765_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold802 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold803 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold804 (.A(_00203_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold805 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold806 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold807 (.A(_01170_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold808 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold809 (.A(_00699_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold810 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold811 (.A(_00217_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold812 (.A(\i_exotiny._0018_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold813 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold814 (.A(_00410_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold815 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold816 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold817 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold818 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold819 (.A(_00779_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold820 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold821 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold822 (.A(_00536_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold823 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold824 (.A(_00456_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold825 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold826 (.A(_00899_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold827 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold828 (.A(_00997_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold829 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold830 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold831 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold832 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold833 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold834 (.A(_00920_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold835 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold836 (.A(_01016_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold837 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold838 (.A(_00312_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold839 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold840 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold841 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold842 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold843 (.A(_00197_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold844 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold845 (.A(_00377_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold846 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold847 (.A(_00438_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold848 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold849 (.A(_00144_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold850 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold851 (.A(_00732_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold852 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold853 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold854 (.A(_01290_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold855 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold856 (.A(_00311_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold857 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold858 (.A(_01337_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold859 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold860 (.A(_01145_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold861 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold862 (.A(_00707_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold863 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold864 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold865 (.A(_00292_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold866 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold867 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold868 (.A(_00851_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold869 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold870 (.A(_01258_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold871 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold872 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold873 (.A(_00239_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold874 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold875 (.A(_00602_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold876 (.A(\i_exotiny._0041_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold877 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold878 (.A(_01295_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold879 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold880 (.A(_01146_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold881 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold882 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold883 (.A(_00306_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold884 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold885 (.A(_00915_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold886 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold887 (.A(_00981_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold888 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold889 (.A(_01004_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold890 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold891 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold892 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold893 (.A(\i_exotiny._0029_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold894 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold895 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold896 (.A(_00743_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold897 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold898 (.A(_01205_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold899 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold900 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold901 (.A(_01192_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold902 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold903 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold904 (.A(_00468_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold905 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold906 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold907 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold908 (.A(\i_exotiny._0369_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold909 (.A(\i_exotiny._1611_[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold910 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold911 (.A(_00538_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold912 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold913 (.A(_00325_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold914 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold915 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold916 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold917 (.A(_01244_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold918 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold919 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold920 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold921 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold922 (.A(_01220_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold923 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold924 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold925 (.A(_01279_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold926 (.A(\i_exotiny._0043_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold927 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold928 (.A(_00200_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold929 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold930 (.A(_00280_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold931 (.A(\i_exotiny._0013_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold932 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold933 (.A(_00984_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold934 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold935 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold936 (.A(_00290_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold937 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold938 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold939 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold940 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold941 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold942 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold943 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold944 (.A(_00753_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold945 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold946 (.A(_00173_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold947 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold948 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold949 (.A(_00421_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold950 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold951 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold952 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold953 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold954 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold955 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold956 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold957 (.A(_00709_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold958 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold959 (.A(_01151_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold960 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold961 (.A(_00901_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold962 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold963 (.A(_01003_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold964 (.A(\i_exotiny._0038_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold965 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold966 (.A(_00156_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold967 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold968 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold969 (.A(_00246_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold970 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold971 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold972 (.A(_00270_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold973 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold974 (.A(_00248_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold975 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold976 (.A(\i_exotiny._0034_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold977 (.A(\i_exotiny._0021_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold978 (.A(\i_exotiny._0034_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold979 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold980 (.A(_00820_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold981 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold982 (.A(_01309_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold983 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold984 (.A(_01354_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold985 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold986 (.A(_00172_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold987 (.A(\i_exotiny._0016_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold988 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold989 (.A(_00081_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold990 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold991 (.A(_00122_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold992 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold993 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold994 (.A(_00430_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold995 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold996 (.A(_00155_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold997 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold998 (.A(_00592_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold999 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold1000 (.A(_00454_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold1001 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold1002 (.A(_00900_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold1003 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold1004 (.A(_00815_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold1007 (.A(_01274_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold1009 (.A(_00590_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold1011 (.A(_01253_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\i_exotiny._0042_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold1014 (.A(\i_exotiny._0315_[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold1015 (.A(_01090_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold1018 (.A(_00262_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold1020 (.A(_01011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold1022 (.A(_00710_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold1025 (.A(_00490_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_01264_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold1029 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold1030 (.A(_00708_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold1032 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold1033 (.A(_01142_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold1035 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\i_exotiny._0314_[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold1038 (.A(_00641_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\i_exotiny._0017_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold1040 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold1041 (.A(_00114_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold1042 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold1043 (.A(_01281_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\i_exotiny._0033_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold1048 (.A(_00598_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold1050 (.A(_00567_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold1052 (.A(_00968_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold1056 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold1057 (.A(_00125_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\i_exotiny._0314_[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold1060 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold1063 (.A(_00961_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold1064 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold1066 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold1069 (.A(_00115_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold1074 (.A(_01242_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold1076 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold1077 (.A(_00123_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold1079 (.A(_00522_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold1080 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold1082 (.A(_00751_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold1083 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold1084 (.A(_01326_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold1086 (.A(_00782_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold1087 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold1091 (.A(_01138_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold1094 (.A(_00801_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold1096 (.A(_01315_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold1098 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold1099 (.A(_00754_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold1101 (.A(_00725_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold1103 (.A(_00483_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold1104 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold1105 (.A(_00120_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\i_exotiny._0038_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold1107 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold1109 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold1110 (.A(_00856_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold1111 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold1114 (.A(_00573_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold1117 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold1119 (.A(\i_exotiny._0013_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold1123 (.A(_00461_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold1124 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold1130 (.A(_00918_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold1135 (.A(_00284_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\i_exotiny._0026_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold1139 (.A(_00612_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold1141 (.A(_00843_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold1143 (.A(_00154_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold1150 (.A(_01195_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold1151 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold1153 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\i_exotiny._0013_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold1157 (.A(_00559_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\i_exotiny._0029_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold1160 (.A(_00387_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold1162 (.A(_00744_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold1164 (.A(_01203_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold1166 (.A(_01199_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold1169 (.A(_00499_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\i_exotiny._0369_[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\i_exotiny._1611_[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold1172 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold1174 (.A(_00831_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\i_exotiny._0015_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\i_exotiny._0024_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold1181 (.A(_01261_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\i_exotiny._0030_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\i_exotiny._1160_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\i_exotiny._0042_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold1188 (.A(_00294_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold1190 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold1191 (.A(_01293_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold1193 (.A(_00563_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold1197 (.A(_00343_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold1200 (.A(_00413_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold1202 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold1203 (.A(_00145_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold1204 (.A(\i_exotiny._0043_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold1206 (.A(_00715_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold1208 (.A(_00773_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold1213 (.A(_00832_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold1215 (.A(_00714_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\i_exotiny._0029_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\i_exotiny._0014_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold1218 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold1219 (.A(_00813_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\i_exotiny._0040_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold1224 (.A(_01262_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\i_exotiny._0315_[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold1228 (.A(_00603_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold1231 (.A(_01243_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold1234 (.A(_00232_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold1236 (.A(\i_exotiny._0015_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\i_exotiny._0039_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\i_exotiny._0017_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold1240 (.A(_01359_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold1242 (.A(_00542_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold1245 (.A(_00988_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold1247 (.A(_00833_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\i_exotiny._0027_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold1249 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold1251 (.A(_00793_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\i_exotiny._0015_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_00147_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold1257 (.A(_00962_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold1259 (.A(_01163_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold1260 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold1261 (.A(_00385_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold1262 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold1264 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold1268 (.A(_00588_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold1271 (.A(_01358_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold1273 (.A(_00739_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold1276 (.A(_00317_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold1277 (.A(\i_exotiny._0034_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold1279 (.A(_01135_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold1283 (.A(_00802_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold1284 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold1285 (.A(_00282_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold1286 (.A(\i_exotiny._0315_[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold1287 (.A(_01092_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold1288 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold1289 (.A(_00545_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold1290 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold1291 (.A(_00585_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold1294 (.A(_00140_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\i_exotiny._0031_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold1297 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold1298 (.A(_01302_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold1300 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold1301 (.A(_00314_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold1302 (.A(\i_exotiny._0017_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold1304 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\i_exotiny._0041_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold1312 (.A(_01180_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold1314 (.A(_01336_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\i_exotiny._1612_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold1316 (.A(_00208_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold1318 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold1319 (.A(_01166_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold1320 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold1321 (.A(_00472_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold1325 (.A(_00546_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold1327 (.A(_00594_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\i_exotiny._0314_[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold1329 (.A(_00647_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold1331 (.A(_01233_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold1334 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold1335 (.A(_00344_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold1338 (.A(_00408_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\i_exotiny._0042_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold1346 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold1348 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold1350 (.A(_01206_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold1352 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold1353 (.A(_00411_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold1355 (.A(_01181_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold1357 (.A(_00786_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold1358 (.A(\i_exotiny._0315_[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\i_exotiny._0029_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold1362 (.A(_00362_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold1365 (.A(_00322_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold1366 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold1373 (.A(_00810_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\i_exotiny._0032_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold1377 (.A(_01266_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold1380 (.A(_00437_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold1382 (.A(_00378_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold1384 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\i_exotiny._0028_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold1388 (.A(_00905_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold1390 (.A(_00741_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\i_exotiny._0315_[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold1394 (.A(_01095_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold1399 (.A(_01285_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold1401 (.A(_01265_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold1403 (.A(_00433_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\i_exotiny._0031_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold1406 (.A(_01020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold1407 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold1409 (.A(_03174_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold1410 (.A(_01128_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[9].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold1413 (.A(_00616_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\i_exotiny.core_res_en_n ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold1415 (.A(_01444_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\i_exotiny._0314_[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold1417 (.A(_00643_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold1419 (.A(_00326_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold1421 (.A(_00738_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\i_exotiny._0023_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold1424 (.A(_01343_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold1426 (.A(_01319_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold1431 (.A(_00457_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\i_exotiny._0014_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold1435 (.A(_00480_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold1438 (.A(_00198_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold1440 (.A(_00458_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\i_exotiny._0028_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold1443 (.A(\i_exotiny._0026_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold1445 (.A(_01209_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold1446 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\i_exotiny._0016_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold1449 (.A(_00817_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold1451 (.A(_00319_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold1453 (.A(_00267_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold1455 (.A(\i_exotiny._0018_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold1457 (.A(_00160_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold1459 (.A(_00393_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold1460 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold1462 (.A(_00742_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold1464 (.A(\i_exotiny._0039_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold1466 (.A(_01272_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\i_exotiny._0027_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold1471 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold1473 (.A(_00713_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold1476 (.A(_00310_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold1478 (.A(_00823_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold1479 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\i_exotiny._0369_[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold1481 (.A(\i_exotiny._1611_[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold1483 (.A(_00735_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold1485 (.A(_01152_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold1488 (.A(_00964_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\i_exotiny._0315_[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold1492 (.A(\i_exotiny._0030_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\i_exotiny._0032_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold1494 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[22].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold1498 (.A(_00503_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.genblk7.g_value.r_value [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold1500 (.A(_02106_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold1501 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold1502 (.A(_00550_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold1504 (.A(_00842_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold1506 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold1509 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\i_exotiny._0033_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[20].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold1512 (.A(_01149_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold1513 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\i_exotiny._0040_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\i_exotiny._0035_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold1517 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold1518 (.A(_00525_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[5].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold1520 (.A(_00553_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold1523 (.A(_00254_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold1526 (.A(_00975_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold1528 (.A(_00488_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\i_exotiny._0314_[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold1532 (.A(_00644_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\i_exotiny._1160_[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold1534 (.A(_01062_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold1537 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold1538 (.A(_00837_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold1542 (.A(_00828_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_00109_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold1547 (.A(_00481_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold1549 (.A(_01294_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\i_exotiny._0315_[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[25].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold1554 (.A(_00711_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\i_exotiny._0314_[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold1556 (.A(_00633_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\i_exotiny._1160_[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold1558 (.A(_01061_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[6].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\i_exotiny._1840_[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\i_exotiny._1611_[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\i_exotiny._0314_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\i_exotiny._1465_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[16].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold1567 (.A(_00315_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold1568 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold1569 (.A(_00783_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\i_exotiny._0036_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold1573 (.A(_02387_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold1574 (.A(_00064_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\i_exotiny._0314_[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold1576 (.A(_00642_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[13].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold1579 (.A(_00426_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\i_exotiny._0314_[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold1581 (.A(_00630_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\i_exotiny._0018_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold1585 (.A(\i_exotiny._0038_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold1587 (.A(_00847_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\i_exotiny._1160_[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold1589 (.A(_01063_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold1591 (.A(_00176_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\i_exotiny._0035_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold1593 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold1594 (.A(_01316_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\i_exotiny._1618_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_00814_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold1603 (.A(\i_exotiny._2025_[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\i_exotiny._1902_[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold1606 (.A(_00487_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[26].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[2].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold1611 (.A(_00922_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[24].i_reg.reg_r[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\i_exotiny._0037_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\i_exotiny._0369_[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\i_exotiny._1611_[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold1618 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold1620 (.A(\i_exotiny._0314_[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold1621 (.A(_00640_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold1623 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold1624 (.A(_00296_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\i_exotiny._0032_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold1629 (.A(_00375_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\i_exotiny._0369_[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\i_exotiny._1611_[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\i_exotiny._0027_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold1633 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[17].i_reg.reg_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[4].i_reg.reg_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\i_exotiny._0314_[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold1636 (.A(_00638_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold1638 (.A(_00853_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\i_exotiny._1586_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold1640 (.A(_00696_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[15].i_reg.reg_r[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold1643 (.A(_01499_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[8].i_reg.reg_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold1645 (.A(_01015_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[18].i_reg.reg_r[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold1647 (.A(_01341_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\i_exotiny._0314_[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\i_exotiny._0314_[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold1650 (.A(_00632_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold1653 (.A(_00358_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[7].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold1656 (.A(_00556_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold1659 (.A(_00218_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold1661 (.A(_00193_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\i_exotiny._0314_[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[23].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[19].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold1665 (.A(_01298_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\i_exotiny._0314_[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold1667 (.A(_00628_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[29].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold1669 (.A(_00354_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold1670 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[28].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\i_exotiny._0314_[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold1672 (.A(_00639_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[21].i_reg.reg_r[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\i_exotiny._1616_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold1675 (.A(_00684_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[3].i_reg.reg_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\i_exotiny._0314_[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\i_exotiny._0369_[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\i_exotiny._1611_[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[12].i_reg.reg_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[1].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold1682 (.A(\i_exotiny._0314_[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\i_exotiny._0033_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold1684 (.A(_00014_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold1685 (.A(_00025_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold1687 (.A(_00204_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[27].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold1689 (.A(_00380_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\i_exotiny._0314_[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold1691 (.A(_00635_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[11].i_reg.reg_r[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\i_exotiny._1715_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold1694 (.A(_01494_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold1695 (.A(_00007_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold1697 (.A(\i_exotiny._1489_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\i_exotiny._0023_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\i_exotiny._1160_[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold1700 (.A(_01048_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\i_exotiny.i_wdg_top.o_wb_dat[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold1702 (.A(_00069_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\i_exotiny.i_wb_spi.dat_rx_r[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold1704 (.A(_00959_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[10].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[31].i_reg.reg_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold1707 (.A(_00919_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold1708 (.A(\i_exotiny._1160_[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold1709 (.A(_01058_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\i_exotiny._0315_[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold1711 (.A(_01076_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[30].i_reg.reg_r[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold1713 (.A(_00478_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold1714 (.A(\i_exotiny._1160_[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold1715 (.A(_01053_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold1716 (.A(_00021_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold1717 (.A(_00214_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\i_exotiny._0315_[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold1719 (.A(_01083_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\i_exotiny._0315_[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold1721 (.A(_01084_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\i_exotiny._0315_[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold1723 (.A(_01088_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\i_exotiny._2025_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\i_exotiny._1902_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\i_exotiny.i_wdg_top.o_wb_dat[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold1727 (.A(_00067_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\i_exotiny._0315_[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold1729 (.A(\i_exotiny.i_wb_spi.dat_rx_r[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold1730 (.A(_00932_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\i_exotiny._1160_[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold1732 (.A(\i_exotiny._1615_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold1733 (.A(_00212_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold1734 (.A(\i_exotiny._2025_[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\i_exotiny._1902_[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\i_exotiny._1617_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold1737 (.A(_00682_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\i_exotiny._1160_[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold1739 (.A(_01055_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold1741 (.A(_00024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold1742 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\i_exotiny._0315_[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold1744 (.A(\i_exotiny.i_rstctl.sys_res_n ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\i_exotiny._1616_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold1746 (.A(_00685_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\i_exotiny.i_wb_spi.dat_rx_r[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold1748 (.A(_00931_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\i_exotiny.i_wb_spi.dat_rx_r[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold1750 (.A(_00930_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold1752 (.A(_03171_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\i_exotiny._0079_[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold1754 (.A(_01069_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\i_exotiny.i_wb_spi.dat_rx_r[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold1756 (.A(_00958_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\i_exotiny._0369_[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\i_exotiny._1611_[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold1759 (.A(\i_exotiny.i_rstctl.cnt[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\i_exotiny.i_wb_spi.dat_rx_r[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold1761 (.A(_00951_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\i_exotiny.i_wb_spi.dat_rx_r[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold1763 (.A(_00929_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold1765 (.A(_00618_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1[14].i_reg.reg_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\i_exotiny._0369_[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\i_exotiny._1611_[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\i_exotiny._0369_[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\i_exotiny._1611_[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold1771 (.A(\i_exotiny._1160_[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold1772 (.A(_01057_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\i_exotiny.i_wb_spi.dat_rx_r[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\i_exotiny._0369_[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\i_exotiny._1611_[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\i_exotiny._0314_[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold1777 (.A(_00629_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\i_exotiny._0314_[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold1779 (.A(\i_exotiny._1956_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold1781 (.A(_03168_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\i_exotiny._1160_[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\i_exotiny._0314_[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\i_exotiny._0315_[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold1786 (.A(_01085_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\i_exotiny._1616_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold1788 (.A(_00686_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\i_exotiny.i_wb_spi.dat_rx_r[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold1790 (.A(_00955_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\i_exotiny._2025_[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\i_exotiny._1902_[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\i_exotiny._1616_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold1794 (.A(_00687_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\i_exotiny._1615_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold1796 (.A(\i_exotiny.i_wb_spi.dat_rx_r[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold1798 (.A(\i_exotiny._0315_[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\i_exotiny._0315_[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold1801 (.A(_03160_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold1802 (.A(_01119_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\i_exotiny._1614_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold1804 (.A(_00678_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\i_exotiny._6090_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold1806 (.A(_00660_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\i_exotiny.i_wb_spi.state_r[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold1808 (.A(_00859_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\i_exotiny._1160_[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\i_exotiny.i_wb_spi.dat_rx_r[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold1812 (.A(_00952_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\i_exotiny.i_wb_spi.state_r[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\i_exotiny._0369_[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\i_exotiny._0369_[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\i_exotiny.i_wb_spi.dat_rx_r[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold1818 (.A(_00948_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\i_exotiny.i_wb_spi.dat_rx_r[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\i_exotiny._0369_[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold1821 (.A(_02575_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold1823 (.A(_03178_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\i_exotiny._1793_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold1825 (.A(_01547_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold1826 (.A(_00010_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold1827 (.A(\i_exotiny.i_wb_spi.dat_rx_r[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\i_exotiny.i_wb_spi.dat_rx_r[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\i_exotiny.i_wb_regs.spi_auto_cs_o ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\i_exotiny._6090_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\i_exotiny.i_rstctl.cnt[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\i_exotiny.i_wb_spi.dat_rx_r[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold1833 (.A(_00954_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\i_exotiny._0315_[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold1835 (.A(_01086_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\i_exotiny.i_wb_spi.dat_rx_r[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold1837 (.A(_00953_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\i_exotiny._0315_[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\i_exotiny.i_wdg_top.o_wb_dat[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold1840 (.A(_00068_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\i_exotiny._1619_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold1842 (.A(_00688_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\i_exotiny._0315_[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold1845 (.A(\i_exotiny._1619_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold1846 (.A(_00690_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\i_exotiny._0014_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\i_exotiny._0369_[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\i_exotiny._1611_[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold1851 (.A(_02248_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\i_exotiny._1489_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\i_exotiny._1617_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\i_exotiny.i_rstctl.cnt[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold1855 (.A(_02903_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold1856 (.A(_02913_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\i_exotiny._0590_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold1858 (.A(_01028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\i_exotiny._1160_[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold1860 (.A(\i_exotiny._1619_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\i_exotiny._0327_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold1862 (.A(_02597_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold1864 (.A(_01025_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\i_exotiny._0315_[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold1866 (.A(_01077_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\i_exotiny._1311_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold1868 (.A(_01508_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold1869 (.A(_00005_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\i_exotiny._1617_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold1871 (.A(_02826_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\i_exotiny.i_wb_qspi_mem.cnt_r[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold1873 (.A(_03152_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold1874 (.A(_01114_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\i_exotiny._1711_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\i_exotiny.i_wb_spi.cnt_hbit_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold1877 (.A(_00060_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\i_exotiny._1623_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\i_exotiny._0315_[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\i_exotiny._1711_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\i_exotiny.i_wdg_top.o_wb_dat[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold1882 (.A(_02407_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold1883 (.A(_00074_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\i_exotiny._1614_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\i_exotiny._1160_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold1886 (.A(\i_exotiny.i_wb_qspi_mem.cnt_r[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\i_exotiny.i_wdg_top.o_wb_dat[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold1888 (.A(_02405_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold1889 (.A(_00073_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\i_exotiny._1617_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold1891 (.A(_00680_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\i_exotiny._6090_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold1893 (.A(_00662_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\i_exotiny.i_wb_regs.spi_size_o[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold1896 (.A(_03177_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\i_exotiny._1725_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold1898 (.A(_01113_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\i_exotiny._0571_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\i_exotiny.i_wb_spi.cnt_presc_r[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\i_exotiny._0369_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data [0]),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold1904 (.A(_00658_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\i_exotiny._1652_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\i_exotiny.i_wb_regs.spi_size_o[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold1907 (.A(_02819_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\i_exotiny.i_wdg_top.o_wb_dat[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold1909 (.A(_00066_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\i_exotiny._0369_[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\i_exotiny._1611_[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold1912 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold1913 (.A(_01033_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\i_exotiny.gpo[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold1915 (.A(_02958_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold1916 (.A(_00926_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\i_exotiny.gpo[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold1918 (.A(_02959_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold1919 (.A(_00927_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\i_exotiny._1619_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold1921 (.A(_00691_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\i_exotiny._0369_[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\i_exotiny._1611_[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\i_exotiny.i_wdg_top.o_wb_dat[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold1925 (.A(_02403_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold1926 (.A(_00072_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold1927 (.A(\i_exotiny._1309_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold1928 (.A(_00009_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold1929 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold1931 (.A(_00619_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\i_exotiny._0369_[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold1933 (.A(_00513_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\i_exotiny._0550_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\i_exotiny._0315_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\i_exotiny.i_rstctl.cnt[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\i_exotiny._0369_[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold1938 (.A(_00509_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold1939 (.A(\i_exotiny.i_rstctl.cnt[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold1940 (.A(\i_exotiny._0601_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\i_exotiny._0369_[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold1942 (.A(_01026_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold1943 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold1944 (.A(_03011_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\i_exotiny.gpo[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold1946 (.A(_02957_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold1947 (.A(_00925_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold1948 (.A(\i_exotiny.i_wb_qspi_mem.crm_r ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold1949 (.A(_02605_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\i_exotiny.i_wb_spi.dat_rx_r[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\i_exotiny._0369_[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold1952 (.A(_00512_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\i_exotiny.i_wdg_top.do_cnt ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold1954 (.A(_02072_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\i_exotiny._2055_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold1957 (.A(\i_exotiny._0315_[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\i_exotiny.i_wdg_top.o_wb_dat[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold1959 (.A(_00070_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\i_exotiny._0369_[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\i_exotiny._6090_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold1962 (.A(\i_exotiny._0327_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold1963 (.A(_01437_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\i_exotiny.i_wdg_top.o_wb_dat[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold1965 (.A(_02409_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold1966 (.A(_00075_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold1968 (.A(\i_exotiny.i_wdg_top.o_wb_dat[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold1969 (.A(_02401_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold1970 (.A(_00071_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\i_exotiny._0369_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\i_exotiny._1611_[30] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold1973 (.A(\i_exotiny._0369_[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\i_exotiny._1615_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold1976 (.A(_03020_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\i_exotiny._0077_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\i_exotiny.i_wb_spi.sck_r ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold1979 (.A(_01231_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\i_exotiny._0542_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\i_exotiny._1612_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold1982 (.A(_00668_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\i_exotiny._0077_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\i_exotiny._1618_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\i_exotiny._0077_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\i_exotiny.i_wb_spi.cnt_presc_r[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\i_exotiny._1660_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold1989 (.A(\i_exotiny._1618_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold1990 (.A(\i_exotiny._1618_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\i_exotiny._0077_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold1992 (.A(\i_exotiny._1306_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\i_exotiny._0315_[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold1994 (.A(_02745_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold1995 (.A(\i_exotiny._0315_[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold1996 (.A(_01072_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\i_exotiny._0079_[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\i_exotiny._0079_[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\i_exotiny._0369_[20] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold2002 (.A(_02582_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\i_exotiny._1757_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\i_exotiny._0077_[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\i_exotiny._1737_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\i_exotiny.i_wdg_top.o_wb_dat[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold2009 (.A(\i_exotiny._0079_[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\i_exotiny._0079_[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold2011 (.A(\i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\i_exotiny._1308_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold2014 (.A(\i_exotiny._3871_ ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold2016 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\i_exotiny.i_wdg_top.clk_div_inst.cnt[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net3844));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_1028 (.VDD(VPWR),
    .VSS(VGND));
endmodule
