* NGSPICE file created from heichips25_fazyrv_exotiny.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

.subckt heichips25_fazyrv_exotiny VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
X_05903_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[8\]
+ net2931 net975 _00120_ VPWR VGND sg13g2_mux2_1
XFILLER_95_884 VPWR VGND sg13g2_decap_8
X_06883_ net1128 _02888_ _02889_ _02890_ VPWR VGND sg13g2_nor3_1
XFILLER_27_406 VPWR VGND sg13g2_fill_2
X_05834_ net2891 net2666 net1054 _00106_ VPWR VGND sg13g2_mux2_1
X_08622_ net1774 VGND VPWR _00694_ i_exotiny._1618_\[2\] clknet_leaf_29_clk_regs sg13g2_dfrbpq_2
X_05765_ _02394_ i_exotiny._2034_\[2\] net1127 VPWR VGND sg13g2_nand2_1
XFILLER_70_718 VPWR VGND sg13g2_fill_2
X_08553_ net702 VGND VPWR _00627_ i_exotiny._0077_\[4\] clknet_leaf_160_clk_regs sg13g2_dfrbpq_1
X_08484_ net196 VGND VPWR _00558_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[4\]
+ clknet_leaf_109_clk_regs sg13g2_dfrbpq_1
X_07504_ net3318 net3706 net902 _01087_ VPWR VGND sg13g2_mux2_1
X_04716_ net14 _01473_ _01474_ VPWR VGND sg13g2_nor2_1
X_05696_ net1117 i_exotiny._1924_\[24\] _02343_ VPWR VGND sg13g2_nor2b_1
X_07435_ _03079_ net1148 _03044_ net1209 i_exotiny._1160_\[20\] VPWR VGND sg13g2_a22oi_1
X_04647_ VPWR _01409_ net1935 VGND sg13g2_inv_1
X_08522__158 VPWR VGND net158 sg13g2_tiehi
X_07366_ _03025_ _02992_ _02999_ VPWR VGND sg13g2_nand2_2
X_07297_ net3036 net3059 net909 _01014_ VPWR VGND sg13g2_mux2_1
X_09105_ net1297 VGND VPWR _01160_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[25\]
+ clknet_leaf_143_clk_regs sg13g2_dfrbpq_1
X_06317_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[15\]
+ net2826 net1033 _00454_ VPWR VGND sg13g2_mux2_1
X_06248_ net2180 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[18\]
+ net1038 _00397_ VPWR VGND sg13g2_mux2_1
X_09036_ net1366 VGND VPWR _01094_ i_exotiny._0315_\[24\] clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
XFILLER_105_923 VPWR VGND sg13g2_decap_8
XFILLER_104_411 VPWR VGND sg13g2_decap_8
Xhold340 _00316_ VPWR VGND net2167 sg13g2_dlygate4sd3_1
X_06179_ net2591 net3174 net950 _00341_ VPWR VGND sg13g2_mux2_1
Xhold351 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[31\]
+ VPWR VGND net2178 sg13g2_dlygate4sd3_1
Xhold362 _01340_ VPWR VGND net2189 sg13g2_dlygate4sd3_1
Xhold395 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[17\]
+ VPWR VGND net2222 sg13g2_dlygate4sd3_1
Xhold373 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[24\]
+ VPWR VGND net2200 sg13g2_dlygate4sd3_1
Xhold384 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[17\]
+ VPWR VGND net2211 sg13g2_dlygate4sd3_1
XFILLER_104_488 VPWR VGND sg13g2_decap_8
X_08097__597 VPWR VGND net597 sg13g2_tiehi
XFILLER_58_542 VPWR VGND sg13g2_fill_1
Xfanout875 _02472_ net875 VPWR VGND sg13g2_buf_8
Xhold1040 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[6\]
+ VPWR VGND net2867 sg13g2_dlygate4sd3_1
Xhold1051 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[12\]
+ VPWR VGND net2878 sg13g2_dlygate4sd3_1
Xfanout886 net890 net886 VPWR VGND sg13g2_buf_8
XFILLER_58_564 VPWR VGND sg13g2_fill_2
XFILLER_58_553 VPWR VGND sg13g2_fill_1
Xfanout897 net900 net897 VPWR VGND sg13g2_buf_8
Xhold1073 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[9\]
+ VPWR VGND net2900 sg13g2_dlygate4sd3_1
Xhold1062 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[5\]
+ VPWR VGND net2889 sg13g2_dlygate4sd3_1
Xhold1084 _01326_ VPWR VGND net2911 sg13g2_dlygate4sd3_1
XFILLER_93_69 VPWR VGND sg13g2_fill_1
Xhold1095 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[18\]
+ VPWR VGND net2922 sg13g2_dlygate4sd3_1
XFILLER_42_95 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_157_clk_regs clknet_5_18__leaf_clk_regs clknet_leaf_157_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_5_365 VPWR VGND sg13g2_fill_2
XFILLER_6_899 VPWR VGND sg13g2_decap_8
XFILLER_97_1003 VPWR VGND sg13g2_decap_8
XFILLER_36_225 VPWR VGND sg13g2_fill_2
XFILLER_51_217 VPWR VGND sg13g2_fill_1
X_05550_ _02230_ VPWR i_exotiny._1611_\[27\] VGND _02219_ _02234_ sg13g2_o21ai_1
X_05481_ net1872 net1070 i_exotiny._1611_\[6\] VPWR VGND sg13g2_and2_1
X_08952__1030 VPWR VGND net1450 sg13g2_tiehi
X_07220_ _02971_ net1937 net1087 VPWR VGND sg13g2_nand2_1
X_07151_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[12\]
+ net2652 net1012 _00899_ VPWR VGND sg13g2_mux2_1
XFILLER_66_0 VPWR VGND sg13g2_fill_1
X_06102_ net2933 net888 _02519_ _02521_ VPWR VGND sg13g2_mux2_1
X_07082_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[10\]
+ net3364 net916 _00837_ VPWR VGND sg13g2_mux2_1
X_06033_ net3485 i_exotiny._0025_\[1\] net963 _00218_ VPWR VGND sg13g2_mux2_1
XFILLER_102_937 VPWR VGND sg13g2_decap_8
XFILLER_99_486 VPWR VGND sg13g2_decap_8
XFILLER_101_436 VPWR VGND sg13g2_decap_8
X_07984_ net125 VGND VPWR net3506 i_exotiny._0369_\[23\] clknet_leaf_165_clk_regs
+ sg13g2_dfrbpq_2
X_06935_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[15\]
+ net3041 net927 _00714_ VPWR VGND sg13g2_mux2_1
X_06866_ VGND VPWR i_exotiny._1619_\[3\] net1134 _02876_ _02875_ sg13g2_a21oi_1
X_05817_ net2750 net2321 net1056 _00089_ VPWR VGND sg13g2_mux2_1
X_08605_ net1791 VGND VPWR _00677_ i_exotiny._1614_\[1\] clknet_leaf_24_clk_regs sg13g2_dfrbpq_2
X_06797_ _02817_ VPWR _02818_ VGND i_exotiny._0369_\[16\] net1191 sg13g2_o21ai_1
X_08168__510 VPWR VGND net510 sg13g2_tiehi
X_05748_ net3606 _01584_ _02383_ VPWR VGND sg13g2_and2_1
X_08536_ net144 VGND VPWR net2618 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[24\]
+ clknet_leaf_176_clk_regs sg13g2_dfrbpq_1
X_05679_ net1916 net1062 _02330_ VPWR VGND sg13g2_nor2_1
XFILLER_24_987 VPWR VGND sg13g2_fill_1
X_08467_ net213 VGND VPWR _00541_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[19\]
+ clknet_leaf_158_clk_regs sg13g2_dfrbpq_1
X_08398_ net538 VGND VPWR net3619 i_exotiny.i_wb_spi.cnt_presc_r\[4\] clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_1
X_07418_ net1082 _03064_ _03065_ _03066_ VPWR VGND sg13g2_nor3_1
X_08598__1378 VPWR VGND net1798 sg13g2_tiehi
XFILLER_7_619 VPWR VGND sg13g2_fill_2
X_08772__1216 VPWR VGND net1636 sg13g2_tiehi
X_07349_ net3771 VPWR _01034_ VGND net1079 _03010_ sg13g2_o21ai_1
XFILLER_6_129 VPWR VGND sg13g2_fill_1
XFILLER_105_720 VPWR VGND sg13g2_decap_8
X_09019_ net1383 VGND VPWR net3693 i_exotiny._0315_\[7\] clknet_leaf_13_clk_regs sg13g2_dfrbpq_2
Xhold170 _01042_ VPWR VGND net1997 sg13g2_dlygate4sd3_1
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_3_858 VPWR VGND sg13g2_decap_8
XFILLER_2_357 VPWR VGND sg13g2_fill_2
XFILLER_105_797 VPWR VGND sg13g2_decap_8
Xhold181 i_exotiny._0314_\[25\] VPWR VGND net2008 sg13g2_dlygate4sd3_1
Xhold192 _00236_ VPWR VGND net2019 sg13g2_dlygate4sd3_1
XFILLER_104_285 VPWR VGND sg13g2_decap_8
XFILLER_92_128 VPWR VGND sg13g2_fill_2
XFILLER_37_84 VPWR VGND sg13g2_fill_1
XFILLER_46_567 VPWR VGND sg13g2_fill_2
XFILLER_73_375 VPWR VGND sg13g2_fill_1
XFILLER_105_1007 VPWR VGND sg13g2_decap_8
X_08505__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_14_475 VPWR VGND sg13g2_fill_2
XFILLER_30_968 VPWR VGND sg13g2_fill_1
X_08748__1240 VPWR VGND net1660 sg13g2_tiehi
XFILLER_6_685 VPWR VGND sg13g2_fill_2
XFILLER_97_968 VPWR VGND sg13g2_decap_8
XFILLER_96_423 VPWR VGND sg13g2_decap_8
Xhold1809 i_exotiny.i_wb_spi.cnt_hbit_r\[1\] VPWR VGND net3636 sg13g2_dlygate4sd3_1
XFILLER_2_880 VPWR VGND sg13g2_decap_8
X_08512__168 VPWR VGND net168 sg13g2_tiehi
X_04981_ _01706_ i_exotiny._6090_\[0\] i_exotiny._6090_\[2\] i_exotiny._6090_\[1\]
+ i_exotiny._6090_\[3\] net1180 _01713_ VPWR VGND sg13g2_mux4_1
Xclkbuf_leaf_54_clk_regs clknet_5_15__leaf_clk_regs clknet_leaf_54_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_65_832 VPWR VGND sg13g2_fill_2
X_06720_ net1173 VPWR _02753_ VGND net3654 net1187 sg13g2_o21ai_1
XFILLER_37_512 VPWR VGND sg13g2_fill_2
XFILLER_49_394 VPWR VGND sg13g2_fill_1
X_06651_ _02689_ _02437_ _02688_ _02692_ VPWR VGND sg13g2_mux2_1
X_05602_ i_exotiny._1956_ _01571_ _02272_ VPWR VGND sg13g2_nor2_1
XFILLER_64_364 VPWR VGND sg13g2_fill_1
XFILLER_52_537 VPWR VGND sg13g2_fill_1
X_06582_ net1199 _02643_ _02644_ _00634_ VPWR VGND sg13g2_nor3_1
X_08321_ net357 VGND VPWR _00402_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[23\]
+ clknet_leaf_73_clk_regs sg13g2_dfrbpq_1
XFILLER_33_751 VPWR VGND sg13g2_fill_2
X_05533_ net1218 _01520_ _02220_ VPWR VGND sg13g2_and2_1
X_08252_ net425 VGND VPWR net2239 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[19\]
+ clknet_leaf_58_clk_regs sg13g2_dfrbpq_1
X_05464_ _02170_ _02140_ i_exotiny._1618_\[3\] _02135_ i_exotiny._1614_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_07203_ VGND VPWR _01411_ net1088 _00936_ _02963_ sg13g2_a21oi_1
X_05395_ _02112_ _02110_ _02111_ VPWR VGND sg13g2_nand2_1
X_08183_ net494 VGND VPWR net2620 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[14\]
+ clknet_leaf_70_clk_regs sg13g2_dfrbpq_1
X_07134_ net1287 net1843 _00884_ VPWR VGND sg13g2_and2_1
XFILLER_106_517 VPWR VGND sg13g2_decap_8
X_07065_ _02937_ net2806 net1014 _00824_ VPWR VGND sg13g2_mux2_1
XFILLER_88_902 VPWR VGND sg13g2_fill_2
X_06016_ _01465_ _01551_ _02126_ _02502_ VPWR VGND sg13g2_nor3_1
XFILLER_102_745 VPWR VGND sg13g2_decap_8
XFILLER_99_283 VPWR VGND sg13g2_decap_8
XFILLER_101_233 VPWR VGND sg13g2_decap_8
XFILLER_88_979 VPWR VGND sg13g2_decap_8
X_07967_ net1178 VGND VPWR net3710 i_exotiny.i_wdg_top.o_wb_dat\[8\] clknet_leaf_48_clk_regs
+ sg13g2_dfrbpq_1
X_06918_ _02485_ _02532_ _02916_ VPWR VGND sg13g2_nor2_2
X_07898_ net44 VGND VPWR net1 i_exotiny.i_rstctl.sys_res_n clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_55_342 VPWR VGND sg13g2_decap_4
X_08826__1162 VPWR VGND net1582 sg13g2_tiehi
Xclkbuf_5_14__f_clk_regs clknet_4_7_0_clk_regs clknet_5_14__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06849_ net3501 net1099 _02862_ VPWR VGND sg13g2_nor2_1
X_08519_ net161 VGND VPWR _00593_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[7\]
+ clknet_leaf_182_clk_regs sg13g2_dfrbpq_1
XFILLER_99_35 VPWR VGND sg13g2_fill_1
XFILLER_87_1013 VPWR VGND sg13g2_decap_8
XFILLER_3_611 VPWR VGND sg13g2_fill_1
XFILLER_105_550 VPWR VGND sg13g2_decap_8
XFILLER_94_927 VPWR VGND sg13g2_decap_8
XFILLER_19_512 VPWR VGND sg13g2_fill_2
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_61_367 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_172_clk_regs clknet_5_5__leaf_clk_regs clknet_leaf_172_clk_regs VPWR
+ VGND sg13g2_buf_8
Xclkbuf_leaf_101_clk_regs clknet_5_23__leaf_clk_regs clknet_leaf_101_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_14_294 VPWR VGND sg13g2_fill_1
XFILLER_7_961 VPWR VGND sg13g2_decap_8
X_05180_ _01900_ VPWR _01908_ VGND _01904_ _01906_ sg13g2_o21ai_1
Xhold917 _01244_ VPWR VGND net2744 sg13g2_dlygate4sd3_1
X_08258__419 VPWR VGND net419 sg13g2_tiehi
Xhold928 _00200_ VPWR VGND net2755 sg13g2_dlygate4sd3_1
Xhold906 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[26\]
+ VPWR VGND net2733 sg13g2_dlygate4sd3_1
X_08158__520 VPWR VGND net520 sg13g2_tiehi
Xhold939 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[10\]
+ VPWR VGND net2766 sg13g2_dlygate4sd3_1
XFILLER_9_1002 VPWR VGND sg13g2_decap_8
X_08870_ net1532 VGND VPWR _00928_ i_exotiny.i_wb_spi.dat_rx_r\[0\] clknet_leaf_29_clk_regs
+ sg13g2_dfrbpq_1
Xhold1606 _00487_ VPWR VGND net3433 sg13g2_dlygate4sd3_1
X_07821_ net2497 _03221_ net891 _01296_ VPWR VGND sg13g2_mux2_1
Xhold1617 i_exotiny._1611_\[22\] VPWR VGND net3444 sg13g2_dlygate4sd3_1
Xhold1639 i_exotiny._1586_ VPWR VGND net3466 sg13g2_dlygate4sd3_1
Xhold1628 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[28\]
+ VPWR VGND net3455 sg13g2_dlygate4sd3_1
X_07752_ net3224 net3157 net991 _01237_ VPWR VGND sg13g2_mux2_1
X_04964_ _01696_ _01424_ _01436_ VPWR VGND sg13g2_xnor2_1
XFILLER_53_813 VPWR VGND sg13g2_fill_1
X_04895_ net1258 net1260 net1222 _01627_ VGND VPWR _01616_ sg13g2_nor4_2
X_07683_ net3181 net2499 net1001 _01185_ VPWR VGND sg13g2_mux2_1
X_06703_ VPWR VGND _01366_ _02738_ _02719_ _01392_ _00661_ net1068 sg13g2_a221oi_1
X_06634_ net2038 net1159 _02679_ VPWR VGND sg13g2_nor2_1
X_08165__513 VPWR VGND net513 sg13g2_tiehi
X_08304_ net374 VGND VPWR net3088 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[6\]
+ clknet_leaf_72_clk_regs sg13g2_dfrbpq_1
X_06565_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[1\].i_hadd.a_i
+ net1160 _02633_ VPWR VGND sg13g2_nor2_1
XFILLER_100_58 VPWR VGND sg13g2_fill_2
X_06496_ net2363 net2999 net1023 _00577_ VPWR VGND sg13g2_mux2_1
X_09284_ net53 VGND VPWR _01339_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[10\]
+ clknet_leaf_170_clk_regs sg13g2_dfrbpq_1
X_05516_ net1277 i_exotiny._0315_\[11\] _02207_ VPWR VGND sg13g2_nor2b_1
X_08235_ net442 VGND VPWR net2167 i_exotiny._0028_\[2\] clknet_leaf_49_clk_regs sg13g2_dfrbpq_2
X_05447_ VGND VPWR i_exotiny._1615_\[1\] _02136_ _02155_ _02137_ sg13g2_a21oi_1
X_05378_ _02100_ _02099_ _02094_ VPWR VGND sg13g2_nand2b_1
X_08166_ net512 VGND VPWR _00247_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[30\]
+ clknet_leaf_132_clk_regs sg13g2_dfrbpq_1
XFILLER_106_314 VPWR VGND sg13g2_decap_8
X_07117_ net1288 net1846 _00867_ VPWR VGND sg13g2_and2_1
X_08097_ net597 VGND VPWR net2208 i_exotiny._0013_\[2\] clknet_leaf_122_clk_regs sg13g2_dfrbpq_2
X_07048_ net3045 net3194 net1017 _00809_ VPWR VGND sg13g2_mux2_1
XFILLER_88_776 VPWR VGND sg13g2_fill_2
XFILLER_87_253 VPWR VGND sg13g2_fill_2
X_08999_ net1403 VGND VPWR net3599 i_exotiny._1160_\[20\] clknet_leaf_18_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_47_117 VPWR VGND sg13g2_fill_2
XFILLER_71_621 VPWR VGND sg13g2_fill_1
X_07988__129 VPWR VGND net129 sg13g2_tiehi
XFILLER_43_356 VPWR VGND sg13g2_fill_2
XFILLER_43_367 VPWR VGND sg13g2_fill_1
X_08502__178 VPWR VGND net178 sg13g2_tiehi
XFILLER_11_286 VPWR VGND sg13g2_fill_2
XFILLER_7_246 VPWR VGND sg13g2_fill_1
XFILLER_4_953 VPWR VGND sg13g2_decap_8
XFILLER_106_881 VPWR VGND sg13g2_decap_8
XFILLER_79_776 VPWR VGND sg13g2_fill_1
Xfanout1231 net1232 net1231 VPWR VGND sg13g2_buf_8
Xfanout1220 net1221 net1220 VPWR VGND sg13g2_buf_8
X_08698__1290 VPWR VGND net1710 sg13g2_tiehi
Xfanout1264 net3815 net1264 VPWR VGND sg13g2_buf_8
Xfanout1253 net1254 net1253 VPWR VGND sg13g2_buf_8
Xfanout1242 i_exotiny._0571_ net1242 VPWR VGND sg13g2_buf_8
Xfanout1286 net1287 net1286 VPWR VGND sg13g2_buf_2
Xfanout1275 net1278 net1275 VPWR VGND sg13g2_buf_8
XFILLER_93_289 VPWR VGND sg13g2_decap_8
XFILLER_75_81 VPWR VGND sg13g2_fill_1
XFILLER_53_109 VPWR VGND sg13g2_fill_2
XFILLER_35_813 VPWR VGND sg13g2_fill_2
X_04680_ _01441_ net1266 _01440_ VPWR VGND sg13g2_nand2_1
X_08593__1383 VPWR VGND net1803 sg13g2_tiehi
XFILLER_90_996 VPWR VGND sg13g2_decap_8
X_06350_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[9\]
+ net3261 net1028 _00480_ VPWR VGND sg13g2_mux2_1
X_06281_ net2797 net2832 net940 _00424_ VPWR VGND sg13g2_mux2_1
X_05301_ _02027_ _01654_ i_exotiny._0020_\[0\] _01618_ i_exotiny._0031_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_08020_ net674 VGND VPWR net2544 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[21\]
+ clknet_leaf_67_clk_regs sg13g2_dfrbpq_1
X_05232_ _01960_ _01624_ i_exotiny._0040_\[1\] _01615_ i_exotiny._0021_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold703 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[10\]
+ VPWR VGND net2530 sg13g2_dlygate4sd3_1
Xhold725 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[9\]
+ VPWR VGND net2552 sg13g2_dlygate4sd3_1
Xhold714 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[9\]
+ VPWR VGND net2541 sg13g2_dlygate4sd3_1
Xhold736 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[14\]
+ VPWR VGND net2563 sg13g2_dlygate4sd3_1
X_05163_ _01887_ _01892_ _01893_ VPWR VGND sg13g2_nor2_1
XFILLER_104_818 VPWR VGND sg13g2_decap_8
Xhold747 _00816_ VPWR VGND net2574 sg13g2_dlygate4sd3_1
Xhold758 _00998_ VPWR VGND net2585 sg13g2_dlygate4sd3_1
X_05094_ VGND VPWR _01824_ _01825_ _01820_ _01601_ sg13g2_a21oi_2
Xhold769 _00189_ VPWR VGND net2596 sg13g2_dlygate4sd3_1
XFILLER_103_339 VPWR VGND sg13g2_decap_8
XFILLER_69_220 VPWR VGND sg13g2_fill_1
X_08922_ net1480 VGND VPWR _00980_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[20\]
+ clknet_leaf_64_clk_regs sg13g2_dfrbpq_1
Xhold1403 _00433_ VPWR VGND net3230 sg13g2_dlygate4sd3_1
Xhold1414 i_exotiny.core_res_en_n VPWR VGND net3241 sg13g2_dlygate4sd3_1
X_08853_ net1553 VGND VPWR _00911_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[20\]
+ clknet_leaf_185_clk_regs sg13g2_dfrbpq_1
Xhold1425 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[26\]
+ VPWR VGND net3252 sg13g2_dlygate4sd3_1
Xhold1458 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[18\]
+ VPWR VGND net3285 sg13g2_dlygate4sd3_1
Xhold1447 i_exotiny._0016_\[2\] VPWR VGND net3274 sg13g2_dlygate4sd3_1
X_05996_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[22\]
+ net3264 net1048 _00198_ VPWR VGND sg13g2_mux2_1
Xhold1436 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[7\]
+ VPWR VGND net3263 sg13g2_dlygate4sd3_1
X_07804_ net3218 net2862 net892 _01283_ VPWR VGND sg13g2_mux2_1
X_08784_ net1624 VGND VPWR net3331 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[15\]
+ clknet_leaf_164_clk_regs sg13g2_dfrbpq_1
Xhold1469 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[18\]
+ VPWR VGND net3296 sg13g2_dlygate4sd3_1
X_07735_ net2613 net876 _03199_ _03203_ VPWR VGND sg13g2_mux2_1
X_04947_ VGND VPWR net1245 net1224 _01679_ net1248 sg13g2_a21oi_1
X_09201__780 VPWR VGND net780 sg13g2_tiehi
XFILLER_66_993 VPWR VGND sg13g2_fill_2
XFILLER_53_654 VPWR VGND sg13g2_fill_2
X_07666_ net3319 net2535 net999 _01168_ VPWR VGND sg13g2_mux2_1
XFILLER_25_345 VPWR VGND sg13g2_fill_2
X_04878_ _01610_ net1254 _01421_ VPWR VGND sg13g2_nand2_1
X_07597_ VGND VPWR i_exotiny.i_wdg_top.clk_div_inst.cnt\[9\] _03166_ _03169_ net1877
+ sg13g2_a21oi_1
X_06617_ net3610 net1155 _02668_ VPWR VGND sg13g2_nor2_1
X_06548_ i_exotiny._0369_\[8\] net1213 _02626_ VPWR VGND sg13g2_and2_1
X_09267_ net93 VGND VPWR _01322_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[25\]
+ clknet_leaf_127_clk_regs sg13g2_dfrbpq_1
X_06479_ net2530 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[6\]
+ net1027 _00560_ VPWR VGND sg13g2_mux2_1
X_08218_ net459 VGND VPWR _00299_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[17\]
+ clknet_leaf_153_clk_regs sg13g2_dfrbpq_1
X_09198_ net783 VGND VPWR net2838 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[20\]
+ clknet_leaf_77_clk_regs sg13g2_dfrbpq_1
XFILLER_106_111 VPWR VGND sg13g2_decap_8
X_08149_ net529 VGND VPWR _00230_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[13\]
+ clknet_leaf_132_clk_regs sg13g2_dfrbpq_1
XFILLER_1_901 VPWR VGND sg13g2_decap_8
XFILLER_106_188 VPWR VGND sg13g2_decap_8
XFILLER_1_978 VPWR VGND sg13g2_decap_8
XFILLER_103_895 VPWR VGND sg13g2_decap_8
XFILLER_102_350 VPWR VGND sg13g2_decap_8
Xhold41 i_exotiny.i_wb_spi.state_r\[19\] VPWR VGND net1868 sg13g2_dlygate4sd3_1
Xhold30 i_exotiny.i_wb_spi.state_r\[7\] VPWR VGND net1857 sg13g2_dlygate4sd3_1
Xhold63 i_exotiny.i_wdg_top.clk_div_inst.cnt\[12\] VPWR VGND net1890 sg13g2_dlygate4sd3_1
Xhold52 _01125_ VPWR VGND net1879 sg13g2_dlygate4sd3_1
Xhold74 i_exotiny._1924_\[18\] VPWR VGND net1901 sg13g2_dlygate4sd3_1
Xhold1970 _00071_ VPWR VGND net3797 sg13g2_dlygate4sd3_1
Xhold1981 i_exotiny._1612_\[0\] VPWR VGND net3808 sg13g2_dlygate4sd3_1
Xhold96 _00037_ VPWR VGND net1923 sg13g2_dlygate4sd3_1
XFILLER_63_418 VPWR VGND sg13g2_fill_1
XFILLER_28_150 VPWR VGND sg13g2_fill_1
Xhold85 _01064_ VPWR VGND net1912 sg13g2_dlygate4sd3_1
Xhold1992 i_exotiny._1306_ VPWR VGND net3819 sg13g2_dlygate4sd3_1
X_08248__429 VPWR VGND net429 sg13g2_tiehi
X_08148__530 VPWR VGND net530 sg13g2_tiehi
XFILLER_8_544 VPWR VGND sg13g2_fill_1
XFILLER_99_849 VPWR VGND sg13g2_decap_8
XFILLER_98_348 VPWR VGND sg13g2_decap_8
X_08785__1203 VPWR VGND net1623 sg13g2_tiehi
X_08155__523 VPWR VGND net523 sg13g2_tiehi
Xfanout1072 _01581_ net1072 VPWR VGND sg13g2_buf_8
Xfanout1061 net1067 net1061 VPWR VGND sg13g2_buf_8
Xfanout1050 net1052 net1050 VPWR VGND sg13g2_buf_8
X_05850_ _02425_ net1245 _02439_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_448 VPWR VGND sg13g2_fill_2
Xfanout1083 net1084 net1083 VPWR VGND sg13g2_buf_1
Xfanout1094 _02717_ net1094 VPWR VGND sg13g2_buf_8
X_04801_ _01548_ net1270 net1181 VPWR VGND sg13g2_nand2_1
X_05781_ _02405_ net1126 _01374_ net1145 net3714 VPWR VGND sg13g2_a22oi_1
X_07520_ VGND VPWR _01500_ _02453_ _03118_ _03117_ sg13g2_a21oi_1
X_04732_ net1231 net3713 net1230 _01488_ VPWR VGND sg13g2_nand3_1
XFILLER_50_624 VPWR VGND sg13g2_decap_8
X_07451_ _03090_ net1148 _03026_ net1207 net3360 VPWR VGND sg13g2_a22oi_1
X_04663_ _01420_ _01423_ _01424_ VPWR VGND sg13g2_and2_1
XFILLER_50_668 VPWR VGND sg13g2_fill_2
X_07382_ i_exotiny._0369_\[29\] net1213 _03037_ VPWR VGND sg13g2_and2_1
X_06402_ i_exotiny._0315_\[16\] i_exotiny._0314_\[16\] net1271 _02586_ VPWR VGND sg13g2_mux2_1
XFILLER_22_326 VPWR VGND sg13g2_fill_2
X_06333_ net2971 net2719 net1037 _00470_ VPWR VGND sg13g2_mux2_1
X_08162__516 VPWR VGND net516 sg13g2_tiehi
X_09121_ net861 VGND VPWR net2302 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[9\]
+ clknet_leaf_155_clk_regs sg13g2_dfrbpq_1
X_09052_ net1350 VGND VPWR net2300 i_exotiny.i_rstctl.cnt\[2\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_1
X_06264_ i_exotiny._0031_\[3\] net874 _02546_ _02551_ VPWR VGND sg13g2_mux2_1
X_08003_ net692 VGND VPWR net2086 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[4\]
+ clknet_leaf_67_clk_regs sg13g2_dfrbpq_1
X_06195_ net3495 net3510 net946 _00350_ VPWR VGND sg13g2_mux2_1
Xhold500 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[20\]
+ VPWR VGND net2327 sg13g2_dlygate4sd3_1
X_05215_ _01942_ VPWR _01943_ VGND i_exotiny._0036_\[1\] _01755_ sg13g2_o21ai_1
Xhold511 _00199_ VPWR VGND net2338 sg13g2_dlygate4sd3_1
Xhold522 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[27\]
+ VPWR VGND net2349 sg13g2_dlygate4sd3_1
Xhold544 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[5\]
+ VPWR VGND net2371 sg13g2_dlygate4sd3_1
Xhold533 _00830_ VPWR VGND net2360 sg13g2_dlygate4sd3_1
X_05146_ _01876_ _01654_ i_exotiny._0020_\[2\] _01627_ i_exotiny._0028_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold566 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[16\]
+ VPWR VGND net2393 sg13g2_dlygate4sd3_1
Xhold577 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[12\]
+ VPWR VGND net2404 sg13g2_dlygate4sd3_1
Xhold588 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[11\]
+ VPWR VGND net2415 sg13g2_dlygate4sd3_1
Xhold555 _00535_ VPWR VGND net2382 sg13g2_dlygate4sd3_1
XFILLER_106_24 VPWR VGND sg13g2_decap_8
XFILLER_103_136 VPWR VGND sg13g2_decap_8
XFILLER_98_860 VPWR VGND sg13g2_decap_8
Xhold599 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[8\]
+ VPWR VGND net2426 sg13g2_dlygate4sd3_1
X_05077_ _01809_ _01779_ i_exotiny._0020_\[3\] _01766_ i_exotiny._0030_\[3\] VPWR
+ VGND sg13g2_a22oi_1
Xclkbuf_leaf_9_clk_regs clknet_5_8__leaf_clk_regs clknet_leaf_9_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold1200 _00413_ VPWR VGND net3027 sg13g2_dlygate4sd3_1
X_08905_ net1497 VGND VPWR _00963_ i_exotiny._0040_\[3\] clknet_leaf_113_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_100_854 VPWR VGND sg13g2_decap_8
Xhold1222 i_exotiny._0040_\[3\] VPWR VGND net3049 sg13g2_dlygate4sd3_1
X_08836_ net1572 VGND VPWR net2080 i_exotiny._0036_\[3\] clknet_leaf_181_clk_regs
+ sg13g2_dfrbpq_2
Xhold1211 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[17\]
+ VPWR VGND net3038 sg13g2_dlygate4sd3_1
Xhold1233 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[15\]
+ VPWR VGND net3060 sg13g2_dlygate4sd3_1
Xhold1255 _00147_ VPWR VGND net3082 sg13g2_dlygate4sd3_1
Xhold1244 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[28\]
+ VPWR VGND net3071 sg13g2_dlygate4sd3_1
Xhold1266 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[18\]
+ VPWR VGND net3093 sg13g2_dlygate4sd3_1
X_08767_ net1641 VGND VPWR _00825_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[30\]
+ clknet_leaf_71_clk_regs sg13g2_dfrbpq_1
Xhold1299 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[25\]
+ VPWR VGND net3126 sg13g2_dlygate4sd3_1
Xhold1277 i_exotiny._0034_\[1\] VPWR VGND net3104 sg13g2_dlygate4sd3_1
X_08648__1329 VPWR VGND net1749 sg13g2_tiehi
Xhold1288 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[27\]
+ VPWR VGND net3115 sg13g2_dlygate4sd3_1
X_05979_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[5\]
+ net2586 net1051 _00181_ VPWR VGND sg13g2_mux2_1
X_08698_ net1710 VGND VPWR _00756_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[25\]
+ clknet_leaf_111_clk_regs sg13g2_dfrbpq_1
X_07718_ net2568 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[15\]
+ net995 _01214_ VPWR VGND sg13g2_mux2_1
X_07649_ net2130 net3004 net900 _01157_ VPWR VGND sg13g2_mux2_1
XFILLER_80_281 VPWR VGND sg13g2_fill_2
XFILLER_31_64 VPWR VGND sg13g2_fill_2
X_08906__1076 VPWR VGND net1496 sg13g2_tiehi
Xoutput31 net31 uio_out[5] VPWR VGND sg13g2_buf_1
Xoutput20 net20 uio_oe[2] VPWR VGND sg13g2_buf_1
XFILLER_95_307 VPWR VGND sg13g2_decap_8
XFILLER_1_775 VPWR VGND sg13g2_decap_8
XFILLER_49_735 VPWR VGND sg13g2_fill_2
XFILLER_36_418 VPWR VGND sg13g2_fill_2
XFILLER_63_248 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_79_clk_regs clknet_5_26__leaf_clk_regs clknet_leaf_79_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_60_977 VPWR VGND sg13g2_fill_1
XFILLER_9_864 VPWR VGND sg13g2_fill_1
XFILLER_8_363 VPWR VGND sg13g2_fill_1
X_05000_ VPWR VGND i_exotiny._6090_\[2\] _01731_ net1180 net1201 _01732_ _01704_ sg13g2_a221oi_1
XFILLER_4_580 VPWR VGND sg13g2_fill_2
X_06951_ net2897 _02919_ net924 _00728_ VPWR VGND sg13g2_mux2_1
X_05902_ net2895 net3219 net972 _00119_ VPWR VGND sg13g2_mux2_1
XFILLER_79_381 VPWR VGND sg13g2_fill_2
XFILLER_95_863 VPWR VGND sg13g2_decap_8
XFILLER_94_340 VPWR VGND sg13g2_decap_4
X_08621_ net1775 VGND VPWR _00693_ i_exotiny._1618_\[1\] clknet_leaf_31_clk_regs sg13g2_dfrbpq_2
X_06882_ net1172 VPWR _02889_ VGND net3582 net1186 sg13g2_o21ai_1
XFILLER_11_0 VPWR VGND sg13g2_fill_2
X_05833_ net3370 net3468 net1057 _00105_ VPWR VGND sg13g2_mux2_1
X_05764_ net1144 net3553 _02393_ _00067_ VPWR VGND sg13g2_a21o_1
X_08552_ net104 VGND VPWR _00626_ i_exotiny._0077_\[3\] clknet_leaf_19_clk_regs sg13g2_dfrbpq_2
X_08483_ net197 VGND VPWR net2082 i_exotiny._0041_\[3\] clknet_leaf_106_clk_regs sg13g2_dfrbpq_2
X_07503_ i_exotiny._0315_\[20\] net3661 net901 _01086_ VPWR VGND sg13g2_mux2_1
X_04715_ net1251 net1252 i_exotiny._0590_ _01473_ VPWR VGND _01432_ sg13g2_nand4_1
X_05695_ net1920 net1061 _02342_ VPWR VGND sg13g2_nor2_1
X_07434_ _03078_ _03025_ _03076_ VPWR VGND sg13g2_nand2_1
X_04646_ VPWR _01408_ net1967 VGND sg13g2_inv_1
X_07365_ net2044 _02991_ _03024_ VPWR VGND sg13g2_nor2_1
X_07296_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[21\]
+ net2103 net908 _01013_ VPWR VGND sg13g2_mux2_1
X_06316_ net3257 net3478 net1036 _00453_ VPWR VGND sg13g2_mux2_1
X_09104_ net1298 VGND VPWR _01159_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[24\]
+ clknet_leaf_142_clk_regs sg13g2_dfrbpq_1
X_06247_ net2373 net2894 net1041 _00396_ VPWR VGND sg13g2_mux2_1
X_09035_ net1367 VGND VPWR _01093_ i_exotiny._0315_\[23\] clknet_leaf_181_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_105_902 VPWR VGND sg13g2_decap_8
Xhold341 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[6\]
+ VPWR VGND net2168 sg13g2_dlygate4sd3_1
X_06178_ net3398 net3161 net952 _00340_ VPWR VGND sg13g2_mux2_1
Xhold352 _00758_ VPWR VGND net2179 sg13g2_dlygate4sd3_1
Xhold330 _00202_ VPWR VGND net2157 sg13g2_dlygate4sd3_1
XFILLER_7_8 VPWR VGND sg13g2_fill_1
XFILLER_105_979 VPWR VGND sg13g2_decap_8
Xhold396 _00812_ VPWR VGND net2223 sg13g2_dlygate4sd3_1
Xhold374 _00399_ VPWR VGND net2201 sg13g2_dlygate4sd3_1
XFILLER_89_145 VPWR VGND sg13g2_fill_1
X_08238__439 VPWR VGND net439 sg13g2_tiehi
Xhold385 _01342_ VPWR VGND net2212 sg13g2_dlygate4sd3_1
Xhold363 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[27\]
+ VPWR VGND net2190 sg13g2_dlygate4sd3_1
X_05129_ _01859_ _01790_ i_exotiny._0034_\[2\] _01770_ i_exotiny._0025_\[2\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_104_467 VPWR VGND sg13g2_decap_8
Xfanout876 net880 net876 VPWR VGND sg13g2_buf_8
Xhold1041 _00114_ VPWR VGND net2868 sg13g2_dlygate4sd3_1
Xhold1030 _00708_ VPWR VGND net2857 sg13g2_dlygate4sd3_1
Xfanout898 net900 net898 VPWR VGND sg13g2_buf_8
Xfanout887 net889 net887 VPWR VGND sg13g2_buf_8
Xhold1074 _01242_ VPWR VGND net2901 sg13g2_dlygate4sd3_1
X_08819_ net1589 VGND VPWR _00877_ i_exotiny.i_wb_spi.state_r\[18\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
Xhold1052 _00968_ VPWR VGND net2879 sg13g2_dlygate4sd3_1
Xhold1063 _00961_ VPWR VGND net2890 sg13g2_dlygate4sd3_1
Xhold1085 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[19\]
+ VPWR VGND net2912 sg13g2_dlygate4sd3_1
Xhold1096 _01315_ VPWR VGND net2923 sg13g2_dlygate4sd3_1
XFILLER_27_974 VPWR VGND sg13g2_fill_1
XFILLER_41_410 VPWR VGND sg13g2_fill_1
XFILLER_42_999 VPWR VGND sg13g2_fill_2
XFILLER_5_322 VPWR VGND sg13g2_fill_1
XFILLER_6_878 VPWR VGND sg13g2_decap_8
XFILLER_6_889 VPWR VGND sg13g2_fill_1
XFILLER_3_35 VPWR VGND sg13g2_decap_4
XFILLER_1_550 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_126_clk_regs clknet_5_23__leaf_clk_regs clknet_leaf_126_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_49_510 VPWR VGND sg13g2_fill_2
X_08152__526 VPWR VGND net526 sg13g2_tiehi
XFILLER_3_1019 VPWR VGND sg13g2_decap_8
XFILLER_92_899 VPWR VGND sg13g2_fill_2
XFILLER_33_944 VPWR VGND sg13g2_fill_2
XFILLER_60_763 VPWR VGND sg13g2_fill_1
XFILLER_32_465 VPWR VGND sg13g2_fill_2
X_05480_ VGND VPWR net1225 _02181_ _02179_ _02178_ sg13g2_a21oi_2
XFILLER_20_649 VPWR VGND sg13g2_fill_2
X_07150_ net2858 net2079 net1012 _00898_ VPWR VGND sg13g2_mux2_1
X_06101_ net2435 net3169 net959 _00277_ VPWR VGND sg13g2_mux2_1
X_07081_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[9\]
+ net2144 net913 _00836_ VPWR VGND sg13g2_mux2_1
XFILLER_59_0 VPWR VGND sg13g2_fill_2
X_06032_ net2637 i_exotiny._0025_\[0\] net964 _00217_ VPWR VGND sg13g2_mux2_1
XFILLER_102_916 VPWR VGND sg13g2_decap_8
XFILLER_101_415 VPWR VGND sg13g2_decap_8
XFILLER_99_465 VPWR VGND sg13g2_decap_8
X_07983_ net124 VGND VPWR net3738 i_exotiny._0369_\[22\] clknet_leaf_165_clk_regs
+ sg13g2_dfrbpq_2
X_06934_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[14\]
+ net3299 net925 _00713_ VPWR VGND sg13g2_mux2_1
X_08862__1124 VPWR VGND net1544 sg13g2_tiehi
X_06865_ net1129 _02873_ _02874_ _02875_ VPWR VGND sg13g2_nor3_1
X_08604_ net1792 VGND VPWR _00676_ i_exotiny._1614_\[0\] clknet_leaf_24_clk_regs sg13g2_dfrbpq_2
X_05816_ net2282 net2085 net1053 _00088_ VPWR VGND sg13g2_mux2_1
Xclkbuf_5_13__f_clk_regs clknet_4_6_0_clk_regs clknet_5_13__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06796_ VGND VPWR _01416_ net1191 _02817_ _01517_ sg13g2_a21oi_1
X_08535_ net145 VGND VPWR _00609_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[23\]
+ clknet_leaf_182_clk_regs sg13g2_dfrbpq_1
XFILLER_36_760 VPWR VGND sg13g2_fill_1
X_05747_ net1931 VPWR _00061_ VGND net1073 _02382_ sg13g2_o21ai_1
XFILLER_35_292 VPWR VGND sg13g2_fill_2
X_05678_ VGND VPWR net1062 _02329_ _00045_ _02327_ sg13g2_a21oi_1
X_08466_ net214 VGND VPWR _00540_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[18\]
+ clknet_leaf_114_clk_regs sg13g2_dfrbpq_1
X_09301__1115 VPWR VGND net1535 sg13g2_tiehi
XFILLER_24_966 VPWR VGND sg13g2_fill_2
X_08397_ net537 VGND VPWR net3552 i_exotiny.i_wb_spi.cnt_presc_r\[3\] clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_50_262 VPWR VGND sg13g2_fill_2
X_07417_ VGND VPWR i_exotiny._0369_\[16\] net1147 _03065_ _03052_ sg13g2_a21oi_1
X_04629_ net3820 _01391_ VPWR VGND sg13g2_inv_4
X_07348_ _03011_ _03004_ _02626_ net1079 net3770 VPWR VGND sg13g2_a22oi_1
X_07279_ net2438 net2767 net909 _00996_ VPWR VGND sg13g2_mux2_1
XFILLER_3_837 VPWR VGND sg13g2_decap_8
X_09018_ net1384 VGND VPWR net3538 i_exotiny._0315_\[6\] clknet_leaf_5_clk_regs sg13g2_dfrbpq_2
Xhold160 i_exotiny._1924_\[6\] VPWR VGND net1987 sg13g2_dlygate4sd3_1
Xhold171 i_exotiny._1924_\[30\] VPWR VGND net1998 sg13g2_dlygate4sd3_1
XFILLER_105_776 VPWR VGND sg13g2_decap_8
XFILLER_104_264 VPWR VGND sg13g2_decap_8
Xhold182 _00649_ VPWR VGND net2009 sg13g2_dlygate4sd3_1
Xhold193 i_exotiny._1160_\[15\] VPWR VGND net2020 sg13g2_dlygate4sd3_1
XFILLER_59_863 VPWR VGND sg13g2_fill_1
XFILLER_26_292 VPWR VGND sg13g2_fill_1
XFILLER_42_752 VPWR VGND sg13g2_fill_2
XFILLER_52_7 VPWR VGND sg13g2_fill_2
XFILLER_69_616 VPWR VGND sg13g2_fill_2
X_08643__1334 VPWR VGND net1754 sg13g2_tiehi
XFILLER_97_947 VPWR VGND sg13g2_decap_8
X_04980_ net1268 VPWR _01712_ VGND _01425_ _01710_ sg13g2_o21ai_1
XFILLER_37_502 VPWR VGND sg13g2_fill_2
X_06650_ _02691_ net1269 _01466_ VPWR VGND sg13g2_nand2_2
X_05601_ VGND VPWR i_exotiny._1612_\[0\] net1106 _00025_ _02271_ sg13g2_a21oi_1
Xclkbuf_leaf_94_clk_regs clknet_5_28__leaf_clk_regs clknet_leaf_94_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_91_173 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_23_clk_regs clknet_5_12__leaf_clk_regs clknet_leaf_23_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06581_ net3475 net1156 _02644_ VPWR VGND sg13g2_nor2_1
X_08320_ net358 VGND VPWR _00401_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[22\]
+ clknet_leaf_76_clk_regs sg13g2_dfrbpq_1
X_08228__449 VPWR VGND net449 sg13g2_tiehi
X_05532_ net1284 VPWR _02219_ VGND i_exotiny._1711_ _02178_ sg13g2_o21ai_1
X_08251_ net426 VGND VPWR _00332_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[18\]
+ clknet_leaf_49_clk_regs sg13g2_dfrbpq_1
X_05463_ VGND VPWR i_exotiny._1615_\[3\] _02136_ _02169_ _02137_ sg13g2_a21oi_1
X_08901__1081 VPWR VGND net1501 sg13g2_tiehi
X_07202_ net1968 net1088 _02963_ VPWR VGND sg13g2_nor2_1
X_05394_ _01400_ VPWR _02111_ VGND _01398_ _01399_ sg13g2_o21ai_1
X_08182_ net495 VGND VPWR _00263_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[13\]
+ clknet_leaf_111_clk_regs sg13g2_dfrbpq_1
X_07133_ net1286 net1862 _00883_ VPWR VGND sg13g2_and2_1
X_07064_ net3129 net883 _02934_ _02937_ VPWR VGND sg13g2_mux2_1
X_06015_ VGND VPWR net2331 net1106 _00210_ _02501_ sg13g2_a21oi_1
XFILLER_102_713 VPWR VGND sg13g2_fill_2
XFILLER_99_262 VPWR VGND sg13g2_decap_8
XFILLER_102_724 VPWR VGND sg13g2_decap_8
XFILLER_101_212 VPWR VGND sg13g2_decap_8
XFILLER_88_958 VPWR VGND sg13g2_decap_8
X_07966_ net1178 VGND VPWR net3716 i_exotiny.i_wdg_top.o_wb_dat\[7\] clknet_leaf_48_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_101_289 VPWR VGND sg13g2_decap_8
XFILLER_96_991 VPWR VGND sg13g2_decap_8
X_06917_ _00698_ net2571 _02915_ VPWR VGND sg13g2_nand2_1
XFILLER_55_310 VPWR VGND sg13g2_fill_1
X_07897_ net2779 _03233_ net980 _01360_ VPWR VGND sg13g2_mux2_1
XFILLER_82_162 VPWR VGND sg13g2_fill_2
X_06848_ VGND VPWR i_exotiny._1619_\[0\] net1134 _02861_ _02860_ sg13g2_a21oi_1
X_06779_ VGND VPWR _02800_ _02802_ _02803_ net1135 sg13g2_a21oi_1
X_08387__291 VPWR VGND net291 sg13g2_tiehi
X_08518_ net162 VGND VPWR net2825 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[6\]
+ clknet_leaf_183_clk_regs sg13g2_dfrbpq_1
XFILLER_24_741 VPWR VGND sg13g2_fill_1
X_08449_ net231 VGND VPWR _00523_ i_exotiny._0039_\[1\] clknet_leaf_159_clk_regs sg13g2_dfrbpq_2
X_08721__1267 VPWR VGND net1687 sg13g2_tiehi
XFILLER_20_980 VPWR VGND sg13g2_fill_2
XFILLER_3_645 VPWR VGND sg13g2_fill_2
XFILLER_2_177 VPWR VGND sg13g2_fill_2
XFILLER_94_906 VPWR VGND sg13g2_decap_8
XFILLER_78_457 VPWR VGND sg13g2_fill_2
X_08943__1039 VPWR VGND net1459 sg13g2_tiehi
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_94_1018 VPWR VGND sg13g2_decap_8
X_07903__50 VPWR VGND net50 sg13g2_tiehi
XFILLER_42_582 VPWR VGND sg13g2_fill_1
XFILLER_80_93 VPWR VGND sg13g2_fill_1
XFILLER_7_940 VPWR VGND sg13g2_decap_8
Xhold918 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[17\]
+ VPWR VGND net2745 sg13g2_dlygate4sd3_1
Xhold907 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[28\]
+ VPWR VGND net2734 sg13g2_dlygate4sd3_1
X_09281__59 VPWR VGND net59 sg13g2_tiehi
Xclkbuf_leaf_141_clk_regs clknet_5_17__leaf_clk_regs clknet_leaf_141_clk_regs VPWR
+ VGND sg13g2_buf_8
Xhold929 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[30\]
+ VPWR VGND net2756 sg13g2_dlygate4sd3_1
Xhold1607 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[14\]
+ VPWR VGND net3434 sg13g2_dlygate4sd3_1
X_07820_ net3249 net875 _03216_ _03221_ VPWR VGND sg13g2_mux2_1
XFILLER_96_287 VPWR VGND sg13g2_decap_8
X_07751_ net2460 net2964 net988 _01236_ VPWR VGND sg13g2_mux2_1
Xhold1629 _00375_ VPWR VGND net3456 sg13g2_dlygate4sd3_1
X_08919__1063 VPWR VGND net1483 sg13g2_tiehi
Xhold1618 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[14\]
+ VPWR VGND net3445 sg13g2_dlygate4sd3_1
X_06702_ VPWR VGND _02737_ net1137 _02735_ net3553 _02738_ net1181 sg13g2_a221oi_1
X_04963_ _01688_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[1\] _01695_ VPWR
+ VGND sg13g2_xor2_1
X_04894_ net1256 _01616_ _01617_ _01626_ VPWR VGND sg13g2_nor3_2
X_07682_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[17\]
+ net2194 net998 _01184_ VPWR VGND sg13g2_mux2_1
XFILLER_25_516 VPWR VGND sg13g2_fill_2
XFILLER_53_836 VPWR VGND sg13g2_fill_2
X_06633_ net1198 _02677_ _02678_ _00651_ VPWR VGND sg13g2_nor3_1
X_06564_ net1195 _02631_ _02632_ _00628_ VPWR VGND sg13g2_nor3_1
X_08303_ net375 VGND VPWR net2417 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[5\]
+ clknet_leaf_84_clk_regs sg13g2_dfrbpq_1
X_05515_ _02206_ net2061 net1070 VPWR VGND sg13g2_nand2_1
X_06495_ net2659 net3012 net1026 _00576_ VPWR VGND sg13g2_mux2_1
X_09283_ net55 VGND VPWR _01338_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[9\]
+ clknet_leaf_179_clk_regs sg13g2_dfrbpq_1
X_08234_ net443 VGND VPWR net3394 i_exotiny._0028_\[1\] clknet_leaf_56_clk_regs sg13g2_dfrbpq_2
X_05446_ _02154_ i_exotiny._0369_\[5\] net1264 VPWR VGND sg13g2_nand2b_1
XFILLER_21_766 VPWR VGND sg13g2_fill_1
X_05377_ VGND VPWR net1112 _02098_ _02099_ _02096_ sg13g2_a21oi_1
X_08165_ net513 VGND VPWR net2796 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[29\]
+ clknet_leaf_132_clk_regs sg13g2_dfrbpq_1
X_07116_ net1289 net1857 _00866_ VPWR VGND sg13g2_and2_1
X_08096_ net598 VGND VPWR _00177_ i_exotiny._0013_\[1\] clknet_leaf_123_clk_regs sg13g2_dfrbpq_2
X_07047_ net2222 net1828 net1015 _00808_ VPWR VGND sg13g2_mux2_1
XFILLER_102_576 VPWR VGND sg13g2_fill_1
XFILLER_88_799 VPWR VGND sg13g2_fill_1
X_07937__711 VPWR VGND net711 sg13g2_tiehi
X_08998_ net1404 VGND VPWR _01056_ i_exotiny._1160_\[19\] clknet_leaf_162_clk_regs
+ sg13g2_dfrbpq_1
X_08739__1249 VPWR VGND net1669 sg13g2_tiehi
X_07949_ net707 VGND VPWR net1973 i_exotiny.i_wb_spi.cnt_hbit_r\[4\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_28_321 VPWR VGND sg13g2_fill_2
XFILLER_55_184 VPWR VGND sg13g2_fill_1
XFILLER_16_538 VPWR VGND sg13g2_fill_1
XFILLER_18_98 VPWR VGND sg13g2_fill_2
XFILLER_43_313 VPWR VGND sg13g2_fill_2
XFILLER_8_704 VPWR VGND sg13g2_fill_2
XFILLER_7_225 VPWR VGND sg13g2_fill_1
XFILLER_4_932 VPWR VGND sg13g2_decap_8
XFILLER_106_860 VPWR VGND sg13g2_decap_8
X_08257__420 VPWR VGND net420 sg13g2_tiehi
XFILLER_59_50 VPWR VGND sg13g2_fill_1
Xfanout1232 net3732 net1232 VPWR VGND sg13g2_buf_8
X_08218__459 VPWR VGND net459 sg13g2_tiehi
XFILLER_39_608 VPWR VGND sg13g2_fill_1
Xfanout1221 _01395_ net1221 VPWR VGND sg13g2_buf_8
Xfanout1210 net1211 net1210 VPWR VGND sg13g2_buf_8
XFILLER_78_265 VPWR VGND sg13g2_fill_1
Xfanout1265 net3833 net1265 VPWR VGND sg13g2_buf_8
Xfanout1254 net3469 net1254 VPWR VGND sg13g2_buf_8
Xfanout1243 i_exotiny._0601_ net1243 VPWR VGND sg13g2_buf_8
Xfanout1287 net1289 net1287 VPWR VGND sg13g2_buf_2
XFILLER_78_298 VPWR VGND sg13g2_fill_2
XFILLER_47_641 VPWR VGND sg13g2_fill_1
Xfanout1276 net1277 net1276 VPWR VGND sg13g2_buf_8
XFILLER_19_398 VPWR VGND sg13g2_fill_2
XFILLER_46_184 VPWR VGND sg13g2_fill_2
XFILLER_90_975 VPWR VGND sg13g2_decap_8
X_08264__413 VPWR VGND net413 sg13g2_tiehi
XFILLER_22_508 VPWR VGND sg13g2_fill_2
XFILLER_62_699 VPWR VGND sg13g2_fill_2
X_06280_ net2507 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[12\]
+ net942 _00423_ VPWR VGND sg13g2_mux2_1
X_05300_ _02026_ _02025_ _01643_ _01646_ i_exotiny._0017_\[0\] VPWR VGND sg13g2_a22oi_1
X_05231_ _01959_ _01648_ i_exotiny._0033_\[1\] _01647_ i_exotiny._0032_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold726 _00121_ VPWR VGND net2553 sg13g2_dlygate4sd3_1
Xhold704 _00560_ VPWR VGND net2531 sg13g2_dlygate4sd3_1
Xhold715 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[27\]
+ VPWR VGND net2542 sg13g2_dlygate4sd3_1
Xhold737 _00231_ VPWR VGND net2564 sg13g2_dlygate4sd3_1
X_05162_ _01889_ _01890_ _01888_ _01892_ VPWR VGND _01891_ sg13g2_nand4_1
Xhold748 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[31\]
+ VPWR VGND net2575 sg13g2_dlygate4sd3_1
X_05093_ _01461_ _01469_ _01822_ _01823_ _01824_ VPWR VGND sg13g2_or4_1
Xhold759 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[9\]
+ VPWR VGND net2586 sg13g2_dlygate4sd3_1
XFILLER_103_318 VPWR VGND sg13g2_decap_8
X_08921_ net1481 VGND VPWR net2455 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[19\]
+ clknet_leaf_66_clk_regs sg13g2_dfrbpq_1
X_08852_ net1554 VGND VPWR _00910_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[19\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
Xhold1404 i_exotiny._0031_\[2\] VPWR VGND net3231 sg13g2_dlygate4sd3_1
Xhold1415 _01444_ VPWR VGND net3242 sg13g2_dlygate4sd3_1
X_07803_ net2625 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[21\]
+ net894 _01282_ VPWR VGND sg13g2_mux2_1
Xhold1459 _00393_ VPWR VGND net3286 sg13g2_dlygate4sd3_1
Xhold1448 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[26\]
+ VPWR VGND net3275 sg13g2_dlygate4sd3_1
XFILLER_84_224 VPWR VGND sg13g2_fill_2
XFILLER_66_950 VPWR VGND sg13g2_fill_2
Xhold1437 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[26\]
+ VPWR VGND net3264 sg13g2_dlygate4sd3_1
X_08783_ net1625 VGND VPWR _00841_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[14\]
+ clknet_leaf_163_clk_regs sg13g2_dfrbpq_1
Xhold1426 _01319_ VPWR VGND net3253 sg13g2_dlygate4sd3_1
X_05995_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[21\]
+ net2669 net1049 _00197_ VPWR VGND sg13g2_mux2_1
XFILLER_72_419 VPWR VGND sg13g2_fill_2
X_07734_ _03202_ net2379 net994 _01228_ VPWR VGND sg13g2_mux2_1
X_04946_ net1245 _01422_ _01678_ VPWR VGND sg13g2_nor2_1
XFILLER_93_780 VPWR VGND sg13g2_fill_2
XFILLER_77_1024 VPWR VGND sg13g2_decap_4
X_07665_ i_exotiny._0030_\[0\] net2182 net1000 _01167_ VPWR VGND sg13g2_mux2_1
X_06616_ net3402 net1163 _02667_ VPWR VGND sg13g2_nor2_1
X_04877_ _01466_ VPWR _01609_ VGND net1252 _01602_ sg13g2_o21ai_1
X_07596_ net1205 net3608 _01124_ VPWR VGND sg13g2_nor2_1
X_08384__294 VPWR VGND net294 sg13g2_tiehi
X_06547_ i_exotiny._0369_\[7\] net3591 net1210 _00618_ VPWR VGND sg13g2_mux2_1
X_06478_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[9\]
+ net2983 net1025 _00559_ VPWR VGND sg13g2_mux2_1
X_09266_ net97 VGND VPWR _01321_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[24\]
+ clknet_leaf_127_clk_regs sg13g2_dfrbpq_1
X_05429_ _02138_ _02129_ _02136_ VPWR VGND sg13g2_nand2_2
X_08217_ net460 VGND VPWR _00298_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[16\]
+ clknet_leaf_171_clk_regs sg13g2_dfrbpq_1
X_08630__1348 VPWR VGND net1768 sg13g2_tiehi
XFILLER_101_1011 VPWR VGND sg13g2_decap_8
X_09197_ net784 VGND VPWR _01252_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[19\]
+ clknet_leaf_77_clk_regs sg13g2_dfrbpq_1
X_08148_ net530 VGND VPWR _00229_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[12\]
+ clknet_leaf_131_clk_regs sg13g2_dfrbpq_1
X_08079_ net615 VGND VPWR net3284 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[16\]
+ clknet_leaf_92_clk_regs sg13g2_dfrbpq_1
XFILLER_84_1028 VPWR VGND sg13g2_fill_1
XFILLER_84_1017 VPWR VGND sg13g2_decap_8
XFILLER_106_167 VPWR VGND sg13g2_decap_8
XFILLER_96_59 VPWR VGND sg13g2_fill_1
XFILLER_1_957 VPWR VGND sg13g2_decap_8
X_08391__287 VPWR VGND net287 sg13g2_tiehi
XFILLER_103_874 VPWR VGND sg13g2_decap_8
Xhold31 i_exotiny.i_wb_spi.state_r\[11\] VPWR VGND net1858 sg13g2_dlygate4sd3_1
Xhold20 i_exotiny.i_wb_spi.state_r\[9\] VPWR VGND net1847 sg13g2_dlygate4sd3_1
XFILLER_0_467 VPWR VGND sg13g2_fill_1
Xhold42 i_exotiny.i_wb_spi.state_r\[4\] VPWR VGND net1869 sg13g2_dlygate4sd3_1
Xhold53 i_exotiny.i_wdg_top.clk_div_inst.cnt\[16\] VPWR VGND net1880 sg13g2_dlygate4sd3_1
Xhold64 _03172_ VPWR VGND net1891 sg13g2_dlygate4sd3_1
Xhold86 i_exotiny.i_wdg_top.clk_div_inst.cnt\[6\] VPWR VGND net1913 sg13g2_dlygate4sd3_1
Xhold75 _00043_ VPWR VGND net1902 sg13g2_dlygate4sd3_1
Xhold97 i_exotiny._1924_\[27\] VPWR VGND net1924 sg13g2_dlygate4sd3_1
Xhold1971 i_exotiny._0369_\[2\] VPWR VGND net3798 sg13g2_dlygate4sd3_1
Xhold1960 i_exotiny._0369_\[16\] VPWR VGND net3787 sg13g2_dlygate4sd3_1
Xhold1982 _00668_ VPWR VGND net3809 sg13g2_dlygate4sd3_1
Xhold1993 i_exotiny._0315_\[4\] VPWR VGND net3820 sg13g2_dlygate4sd3_1
XFILLER_16_313 VPWR VGND sg13g2_fill_1
XFILLER_43_110 VPWR VGND sg13g2_decap_8
X_08893__1089 VPWR VGND net1509 sg13g2_tiehi
XFILLER_101_91 VPWR VGND sg13g2_fill_2
XFILLER_99_828 VPWR VGND sg13g2_decap_8
XFILLER_98_327 VPWR VGND sg13g2_decap_8
XFILLER_79_552 VPWR VGND sg13g2_fill_1
Xfanout1040 net1042 net1040 VPWR VGND sg13g2_buf_8
Xfanout1073 _01581_ net1073 VPWR VGND sg13g2_buf_1
Xfanout1062 net1063 net1062 VPWR VGND sg13g2_buf_8
Xfanout1051 net1052 net1051 VPWR VGND sg13g2_buf_8
X_05780_ _02404_ i_exotiny._2034_\[7\] net1127 VPWR VGND sg13g2_nand2_1
XFILLER_66_268 VPWR VGND sg13g2_fill_1
X_04800_ _00010_ _01546_ net3652 VPWR VGND sg13g2_nand2_1
Xfanout1095 _02717_ net1095 VPWR VGND sg13g2_buf_1
Xfanout1084 net1085 net1084 VPWR VGND sg13g2_buf_2
XFILLER_82_739 VPWR VGND sg13g2_fill_2
X_04731_ _01487_ net1230 net1231 net3713 VPWR VGND sg13g2_and3_2
X_08680__1308 VPWR VGND net1728 sg13g2_tiehi
XFILLER_62_474 VPWR VGND sg13g2_fill_1
X_04662_ net1242 net1247 _01423_ VPWR VGND sg13g2_nor2_2
X_07450_ _03089_ VPWR _01057_ VGND net1082 _03088_ sg13g2_o21ai_1
X_06401_ _02585_ VPWR _00512_ VGND _02572_ _02584_ sg13g2_o21ai_1
X_07381_ VGND VPWR net1077 _03036_ _01041_ _03034_ sg13g2_a21oi_1
XFILLER_89_0 VPWR VGND sg13g2_fill_1
X_06332_ net2353 net2016 net1035 _00469_ VPWR VGND sg13g2_mux2_1
X_09120_ net862 VGND VPWR _01175_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[8\]
+ clknet_leaf_152_clk_regs sg13g2_dfrbpq_1
X_09051_ net1351 VGND VPWR _01106_ i_exotiny.i_rstctl.cnt\[1\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_2
X_07927__721 VPWR VGND net721 sg13g2_tiehi
X_06263_ _02550_ net3136 net1042 _00409_ VPWR VGND sg13g2_mux2_1
X_08002_ net693 VGND VPWR net2215 i_exotiny._0018_\[3\] clknet_leaf_66_clk_regs sg13g2_dfrbpq_2
X_06194_ net2565 net3337 net948 _00349_ VPWR VGND sg13g2_mux2_1
Xhold501 _01345_ VPWR VGND net2328 sg13g2_dlygate4sd3_1
X_05214_ _01938_ _01941_ _01934_ _01942_ VPWR VGND sg13g2_nand3_1
Xhold512 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[18\]
+ VPWR VGND net2339 sg13g2_dlygate4sd3_1
Xhold534 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[10\]
+ VPWR VGND net2361 sg13g2_dlygate4sd3_1
Xhold523 _01158_ VPWR VGND net2350 sg13g2_dlygate4sd3_1
Xhold545 _01330_ VPWR VGND net2372 sg13g2_dlygate4sd3_1
X_05145_ _01875_ _01641_ i_exotiny._0035_\[2\] _01634_ i_exotiny._0013_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold578 _01241_ VPWR VGND net2405 sg13g2_dlygate4sd3_1
Xhold567 _00807_ VPWR VGND net2394 sg13g2_dlygate4sd3_1
Xhold556 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[28\]
+ VPWR VGND net2383 sg13g2_dlygate4sd3_1
XFILLER_1_209 VPWR VGND sg13g2_fill_2
Xhold589 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[9\]
+ VPWR VGND net2416 sg13g2_dlygate4sd3_1
X_05076_ _01808_ _01778_ i_exotiny._0035_\[3\] _01772_ i_exotiny._0033_\[3\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_106_69 VPWR VGND sg13g2_decap_8
XFILLER_100_800 VPWR VGND sg13g2_fill_1
X_08904_ net1498 VGND VPWR net3084 i_exotiny._0040_\[2\] clknet_leaf_65_clk_regs sg13g2_dfrbpq_2
XFILLER_100_833 VPWR VGND sg13g2_decap_8
Xhold1223 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[29\]
+ VPWR VGND net3050 sg13g2_dlygate4sd3_1
XFILLER_58_758 VPWR VGND sg13g2_fill_1
X_08835_ net1573 VGND VPWR _00893_ i_exotiny._0036_\[2\] clknet_leaf_184_clk_regs
+ sg13g2_dfrbpq_2
Xhold1212 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[9\]
+ VPWR VGND net3039 sg13g2_dlygate4sd3_1
Xhold1234 _00232_ VPWR VGND net3061 sg13g2_dlygate4sd3_1
Xhold1201 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[13\]
+ VPWR VGND net3028 sg13g2_dlygate4sd3_1
X_08766_ net1642 VGND VPWR _00824_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[29\]
+ clknet_leaf_82_clk_regs sg13g2_dfrbpq_1
Xhold1245 _00988_ VPWR VGND net3072 sg13g2_dlygate4sd3_1
X_07934__714 VPWR VGND net714 sg13g2_tiehi
Xhold1256 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[6\]
+ VPWR VGND net3083 sg13g2_dlygate4sd3_1
Xhold1267 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[6\]
+ VPWR VGND net3094 sg13g2_dlygate4sd3_1
XFILLER_66_791 VPWR VGND sg13g2_fill_2
X_05978_ net3417 net3484 net1052 _00180_ VPWR VGND sg13g2_mux2_1
X_07717_ net2422 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[14\]
+ net995 _01213_ VPWR VGND sg13g2_mux2_1
X_08656__1321 VPWR VGND net1741 sg13g2_tiehi
Xhold1278 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[4\]
+ VPWR VGND net3105 sg13g2_dlygate4sd3_1
Xhold1289 _00545_ VPWR VGND net3116 sg13g2_dlygate4sd3_1
X_08697_ net1711 VGND VPWR net2356 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[24\]
+ clknet_leaf_104_clk_regs sg13g2_dfrbpq_1
XFILLER_26_655 VPWR VGND sg13g2_fill_1
X_04929_ _01661_ _01636_ i_exotiny._0019_\[3\] _01627_ i_exotiny._0028_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_08247__430 VPWR VGND net430 sg13g2_tiehi
X_07648_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[21\]
+ net2396 net898 _01156_ VPWR VGND sg13g2_mux2_1
XFILLER_25_154 VPWR VGND sg13g2_fill_2
XFILLER_41_625 VPWR VGND sg13g2_fill_1
X_07579_ _03158_ net3844 net1885 _03154_ VPWR VGND sg13g2_and3_1
XFILLER_90_1010 VPWR VGND sg13g2_decap_8
X_08689__1299 VPWR VGND net1719 sg13g2_tiehi
X_08208__469 VPWR VGND net469 sg13g2_tiehi
X_09249_ net558 VGND VPWR _01304_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[7\]
+ clknet_leaf_131_clk_regs sg13g2_dfrbpq_1
X_08878__1104 VPWR VGND net1524 sg13g2_tiehi
XFILLER_31_54 VPWR VGND sg13g2_fill_1
Xoutput21 net21 uio_oe[3] VPWR VGND sg13g2_buf_1
Xoutput32 net32 uio_out[6] VPWR VGND sg13g2_buf_1
X_08254__423 VPWR VGND net423 sg13g2_tiehi
XFILLER_1_754 VPWR VGND sg13g2_decap_8
XFILLER_49_703 VPWR VGND sg13g2_fill_1
XFILLER_64_728 VPWR VGND sg13g2_fill_2
XFILLER_17_600 VPWR VGND sg13g2_fill_2
Xhold1790 _00955_ VPWR VGND net3617 sg13g2_dlygate4sd3_1
XFILLER_32_614 VPWR VGND sg13g2_fill_1
X_08261__416 VPWR VGND net416 sg13g2_tiehi
XFILLER_99_603 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_48_clk_regs clknet_5_14__leaf_clk_regs clknet_leaf_48_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08439__246 VPWR VGND net246 sg13g2_tiehi
X_08734__1254 VPWR VGND net1674 sg13g2_tiehi
X_06950_ net3187 net882 _02916_ _02919_ VPWR VGND sg13g2_mux2_1
X_05901_ net2867 net2817 net975 _00118_ VPWR VGND sg13g2_mux2_1
X_06881_ net3457 net1189 _02888_ VPWR VGND sg13g2_nor2_1
XFILLER_67_577 VPWR VGND sg13g2_fill_2
Xclkbuf_5_12__f_clk_regs clknet_4_6_0_clk_regs clknet_5_12__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_05832_ net3306 net2948 net1053 _00104_ VPWR VGND sg13g2_mux2_1
XFILLER_27_408 VPWR VGND sg13g2_fill_1
X_08620_ net1776 VGND VPWR _00692_ i_exotiny._1618_\[0\] clknet_leaf_8_clk_regs sg13g2_dfrbpq_2
X_05763_ _01399_ net1144 net1143 _02393_ VPWR VGND sg13g2_nor3_1
X_08551_ net105 VGND VPWR _00625_ i_exotiny._0077_\[2\] clknet_leaf_18_clk_regs sg13g2_dfrbpq_2
X_08956__1026 VPWR VGND net1446 sg13g2_tiehi
X_08482_ net198 VGND VPWR net3483 i_exotiny._0041_\[2\] clknet_leaf_108_clk_regs sg13g2_dfrbpq_2
X_05694_ VGND VPWR net1064 _02340_ _00049_ _02341_ sg13g2_a21oi_1
X_07502_ i_exotiny._0315_\[19\] net3612 net904 _01085_ VPWR VGND sg13g2_mux2_1
XFILLER_35_452 VPWR VGND sg13g2_fill_2
X_04714_ i_exotiny._0590_ net1250 net1252 _01432_ _01472_ VPWR VGND sg13g2_and4_1
X_04645_ VPWR _01407_ net3589 VGND sg13g2_inv_1
XFILLER_50_422 VPWR VGND sg13g2_fill_2
X_07433_ _03025_ _03076_ _03077_ VPWR VGND sg13g2_and2_1
XFILLER_50_455 VPWR VGND sg13g2_decap_4
X_09103_ net1299 VGND VPWR net2350 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[23\]
+ clknet_leaf_144_clk_regs sg13g2_dfrbpq_1
X_08381__297 VPWR VGND net297 sg13g2_tiehi
X_07364_ _03023_ VPWR _01037_ VGND net1079 _03022_ sg13g2_o21ai_1
X_07295_ net2245 net2662 net910 _01012_ VPWR VGND sg13g2_mux2_1
X_06315_ net2650 net2538 net1034 _00452_ VPWR VGND sg13g2_mux2_1
X_06246_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[20\]
+ net2621 net1041 _00395_ VPWR VGND sg13g2_mux2_1
X_08277__401 VPWR VGND net401 sg13g2_tiehi
X_09034_ net1368 VGND VPWR net3114 i_exotiny._0315_\[22\] clknet_leaf_179_clk_regs
+ sg13g2_dfrbpq_1
Xhold320 _00347_ VPWR VGND net2147 sg13g2_dlygate4sd3_1
Xhold353 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[22\]
+ VPWR VGND net2180 sg13g2_dlygate4sd3_1
Xhold342 _00146_ VPWR VGND net2169 sg13g2_dlygate4sd3_1
X_06177_ net2226 net3023 net951 _00339_ VPWR VGND sg13g2_mux2_1
Xhold331 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[21\]
+ VPWR VGND net2158 sg13g2_dlygate4sd3_1
XFILLER_105_958 VPWR VGND sg13g2_decap_8
XFILLER_104_446 VPWR VGND sg13g2_decap_8
Xhold375 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[7\]
+ VPWR VGND net2202 sg13g2_dlygate4sd3_1
Xhold386 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[21\]
+ VPWR VGND net2213 sg13g2_dlygate4sd3_1
Xhold364 _01352_ VPWR VGND net2191 sg13g2_dlygate4sd3_1
X_05128_ _01851_ _01856_ _01847_ _01858_ VPWR VGND _01857_ sg13g2_nand4_1
Xhold397 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[19\]
+ VPWR VGND net2224 sg13g2_dlygate4sd3_1
X_05059_ net1221 _01756_ _01757_ _01791_ VPWR VGND sg13g2_nor3_2
Xhold1020 _01011_ VPWR VGND net2847 sg13g2_dlygate4sd3_1
Xfanout888 net889 net888 VPWR VGND sg13g2_buf_8
XFILLER_58_566 VPWR VGND sg13g2_fill_1
Xhold1031 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[11\]
+ VPWR VGND net2858 sg13g2_dlygate4sd3_1
Xhold1042 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[16\]
+ VPWR VGND net2869 sg13g2_dlygate4sd3_1
Xfanout899 net900 net899 VPWR VGND sg13g2_buf_8
Xfanout877 net879 net877 VPWR VGND sg13g2_buf_8
X_08818_ net1590 VGND VPWR net1860 i_exotiny.i_wb_spi.state_r\[17\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
Xhold1053 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[29\]
+ VPWR VGND net2880 sg13g2_dlygate4sd3_1
Xhold1064 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[30\]
+ VPWR VGND net2891 sg13g2_dlygate4sd3_1
X_08605__1371 VPWR VGND net1791 sg13g2_tiehi
Xhold1075 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[14\]
+ VPWR VGND net2902 sg13g2_dlygate4sd3_1
X_08749_ net1659 VGND VPWR net2394 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[12\]
+ clknet_leaf_81_clk_regs sg13g2_dfrbpq_1
Xhold1097 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[17\]
+ VPWR VGND net2924 sg13g2_dlygate4sd3_1
Xhold1086 _00782_ VPWR VGND net2913 sg13g2_dlygate4sd3_1
X_08812__1176 VPWR VGND net1596 sg13g2_tiehi
XFILLER_41_466 VPWR VGND sg13g2_fill_1
XFILLER_6_857 VPWR VGND sg13g2_decap_8
XFILLER_5_367 VPWR VGND sg13g2_fill_1
XFILLER_3_14 VPWR VGND sg13g2_decap_8
X_07917__731 VPWR VGND net731 sg13g2_tiehi
Xclkbuf_leaf_166_clk_regs clknet_5_4__leaf_clk_regs clknet_leaf_166_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_60_786 VPWR VGND sg13g2_fill_2
X_06100_ net2769 net2756 net958 _00276_ VPWR VGND sg13g2_mux2_1
XFILLER_9_695 VPWR VGND sg13g2_fill_2
XFILLER_8_150 VPWR VGND sg13g2_fill_2
X_07080_ net3335 net3076 net913 _00835_ VPWR VGND sg13g2_mux2_1
X_07924__724 VPWR VGND net724 sg13g2_tiehi
X_06031_ VGND VPWR net1138 _02510_ _02511_ net1165 sg13g2_a21oi_1
XFILLER_99_444 VPWR VGND sg13g2_decap_8
X_08237__440 VPWR VGND net440 sg13g2_tiehi
X_07982_ net123 VGND VPWR net3676 i_exotiny._0369_\[21\] clknet_leaf_14_clk_regs sg13g2_dfrbpq_2
XFILLER_68_820 VPWR VGND sg13g2_fill_1
X_06933_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[13\]
+ net2265 net924 _00712_ VPWR VGND sg13g2_mux2_1
X_08574__56 VPWR VGND net56 sg13g2_tiehi
XFILLER_28_706 VPWR VGND sg13g2_fill_2
X_06864_ net1170 VPWR _02874_ VGND net3616 net1186 sg13g2_o21ai_1
X_06795_ _02816_ net3733 _02745_ VPWR VGND sg13g2_nand2_1
X_05815_ net2540 net2214 net1053 _00087_ VPWR VGND sg13g2_mux2_1
X_08603_ net1793 VGND VPWR _00675_ i_exotiny._1615_\[3\] clknet_leaf_23_clk_regs sg13g2_dfrbpq_2
X_05746_ _02374_ VPWR _02382_ VGND net1118 _02381_ sg13g2_o21ai_1
X_07931__717 VPWR VGND net717 sg13g2_tiehi
X_08534_ net146 VGND VPWR _00608_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[22\]
+ clknet_leaf_184_clk_regs sg13g2_dfrbpq_1
XFILLER_36_783 VPWR VGND sg13g2_fill_1
X_05677_ VGND VPWR i_exotiny._1617_\[3\] net1121 _02329_ _02328_ sg13g2_a21oi_1
X_08465_ net215 VGND VPWR _00539_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[17\]
+ clknet_leaf_163_clk_regs sg13g2_dfrbpq_1
X_08244__433 VPWR VGND net433 sg13g2_tiehi
X_08396_ net536 VGND VPWR i_exotiny._1902_\[2\] i_exotiny.i_wb_spi.cnt_presc_r\[2\]
+ clknet_leaf_32_clk_regs sg13g2_dfrbpq_1
X_04628_ net3762 _01390_ VPWR VGND sg13g2_inv_4
XFILLER_23_499 VPWR VGND sg13g2_fill_2
X_07416_ i_exotiny._1160_\[16\] net1216 _03064_ VPWR VGND sg13g2_nor2_1
X_07347_ _03010_ _03008_ _03009_ net1212 net2044 VPWR VGND sg13g2_a22oi_1
X_07278_ i_exotiny._0042_\[3\] net2202 net911 _00995_ VPWR VGND sg13g2_mux2_1
X_09017_ net1385 VGND VPWR _01075_ i_exotiny._0315_\[5\] clknet_leaf_11_clk_regs sg13g2_dfrbpq_2
X_06229_ VGND VPWR net1139 _02546_ _02547_ net1166 sg13g2_a21oi_1
XFILLER_12_89 VPWR VGND sg13g2_fill_2
XFILLER_3_816 VPWR VGND sg13g2_decap_8
XFILLER_105_755 VPWR VGND sg13g2_decap_8
Xhold161 _00031_ VPWR VGND net1988 sg13g2_dlygate4sd3_1
Xhold150 _00459_ VPWR VGND net1977 sg13g2_dlygate4sd3_1
XFILLER_104_243 VPWR VGND sg13g2_decap_8
Xhold172 _00055_ VPWR VGND net1999 sg13g2_dlygate4sd3_1
XFILLER_2_359 VPWR VGND sg13g2_fill_1
Xhold194 _01052_ VPWR VGND net2021 sg13g2_dlygate4sd3_1
Xhold183 i_exotiny._1160_\[13\] VPWR VGND net2010 sg13g2_dlygate4sd3_1
X_08251__426 VPWR VGND net426 sg13g2_tiehi
XFILLER_101_983 VPWR VGND sg13g2_decap_8
XFILLER_100_493 VPWR VGND sg13g2_decap_8
XFILLER_2_1020 VPWR VGND sg13g2_decap_8
XFILLER_18_227 VPWR VGND sg13g2_fill_2
XFILLER_37_75 VPWR VGND sg13g2_decap_8
X_08429__256 VPWR VGND net256 sg13g2_tiehi
XFILLER_46_569 VPWR VGND sg13g2_fill_1
XFILLER_26_271 VPWR VGND sg13g2_fill_1
X_09278__65 VPWR VGND net65 sg13g2_tiehi
XFILLER_14_477 VPWR VGND sg13g2_fill_1
XFILLER_6_643 VPWR VGND sg13g2_fill_1
XFILLER_6_687 VPWR VGND sg13g2_fill_1
X_08436__249 VPWR VGND net249 sg13g2_tiehi
XFILLER_97_926 VPWR VGND sg13g2_decap_8
XFILLER_78_93 VPWR VGND sg13g2_fill_2
XFILLER_65_834 VPWR VGND sg13g2_fill_1
X_05600_ net3511 net1105 _02271_ VPWR VGND sg13g2_nor2_1
X_08267__411 VPWR VGND net411 sg13g2_tiehi
X_06580_ net3407 net1164 _02643_ VPWR VGND sg13g2_nor2_1
XFILLER_45_591 VPWR VGND sg13g2_fill_2
X_05531_ _02218_ net3749 net1071 VPWR VGND sg13g2_nand2_1
X_08250_ net427 VGND VPWR _00331_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[17\]
+ clknet_leaf_48_clk_regs sg13g2_dfrbpq_1
X_05462_ _02168_ i_exotiny._0369_\[7\] net1264 VPWR VGND sg13g2_nand2b_1
X_07201_ VGND VPWR _01410_ net1091 _00935_ _02962_ sg13g2_a21oi_1
Xclkbuf_leaf_63_clk_regs clknet_5_13__leaf_clk_regs clknet_leaf_63_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08181_ net496 VGND VPWR net2845 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[12\]
+ clknet_leaf_110_clk_regs sg13g2_dfrbpq_1
XFILLER_32_296 VPWR VGND sg13g2_fill_1
X_07132_ net1287 net1845 _00882_ VPWR VGND sg13g2_and2_1
X_05393_ i_exotiny._2034_\[1\] i_exotiny._2034_\[2\] i_exotiny._2034_\[0\] _02110_
+ VPWR VGND sg13g2_nand3_1
XFILLER_71_0 VPWR VGND sg13g2_fill_2
X_07063_ _02936_ net3304 net1013 _00823_ VPWR VGND sg13g2_mux2_1
X_06014_ _00017_ net1106 _02501_ VPWR VGND sg13g2_nor2_1
X_08274__404 VPWR VGND net404 sg13g2_tiehi
XFILLER_99_241 VPWR VGND sg13g2_decap_8
XFILLER_88_915 VPWR VGND sg13g2_fill_1
XFILLER_88_904 VPWR VGND sg13g2_fill_1
XFILLER_0_819 VPWR VGND sg13g2_decap_8
XFILLER_87_458 VPWR VGND sg13g2_fill_2
X_07965_ net1177 VGND VPWR net3753 i_exotiny.i_wdg_top.o_wb_dat\[6\] clknet_leaf_48_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_101_268 VPWR VGND sg13g2_decap_8
XFILLER_96_970 VPWR VGND sg13g2_decap_8
X_06916_ VGND VPWR i_exotiny.core_res_en_n _02907_ _02915_ net1227 sg13g2_a21oi_1
XFILLER_68_672 VPWR VGND sg13g2_fill_1
X_07896_ net2804 net872 _03228_ _03233_ VPWR VGND sg13g2_mux2_1
X_06847_ net1129 _02858_ _02859_ _02860_ VPWR VGND sg13g2_nor3_1
XFILLER_15_208 VPWR VGND sg13g2_fill_1
X_06778_ _02801_ VPWR _02802_ VGND net3749 net1190 sg13g2_o21ai_1
X_08998__984 VPWR VGND net1404 sg13g2_tiehi
X_05729_ i_exotiny._1956_ i_exotiny.i_wb_spi.cnt_hbit_r\[1\] i_exotiny.i_wb_spi.cnt_hbit_r\[2\]
+ net1991 _02367_ VPWR VGND sg13g2_nor4_1
XFILLER_51_550 VPWR VGND sg13g2_decap_4
X_08517_ net163 VGND VPWR _00591_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[5\]
+ clknet_leaf_177_clk_regs sg13g2_dfrbpq_1
XFILLER_36_591 VPWR VGND sg13g2_fill_2
X_08448_ net232 VGND VPWR net2906 i_exotiny._0039_\[0\] clknet_leaf_115_clk_regs sg13g2_dfrbpq_2
XFILLER_23_252 VPWR VGND sg13g2_fill_1
X_08379_ net299 VGND VPWR net2114 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[17\]
+ clknet_leaf_139_clk_regs sg13g2_dfrbpq_1
XFILLER_3_635 VPWR VGND sg13g2_fill_1
XFILLER_105_585 VPWR VGND sg13g2_decap_8
X_08951__1031 VPWR VGND net1451 sg13g2_tiehi
XFILLER_78_447 VPWR VGND sg13g2_fill_1
XFILLER_87_992 VPWR VGND sg13g2_decap_8
XFILLER_48_85 VPWR VGND sg13g2_fill_1
XFILLER_59_694 VPWR VGND sg13g2_fill_1
XFILLER_58_193 VPWR VGND sg13g2_fill_2
XFILLER_100_290 VPWR VGND sg13g2_decap_8
X_07914__734 VPWR VGND net734 sg13g2_tiehi
X_08442__242 VPWR VGND net242 sg13g2_tiehi
XFILLER_15_775 VPWR VGND sg13g2_fill_2
XFILLER_42_561 VPWR VGND sg13g2_fill_2
X_08227__450 VPWR VGND net450 sg13g2_tiehi
XFILLER_11_981 VPWR VGND sg13g2_decap_8
Xhold919 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[21\]
+ VPWR VGND net2746 sg13g2_dlygate4sd3_1
Xhold908 i_exotiny._0369_\[1\] VPWR VGND net2735 sg13g2_dlygate4sd3_1
X_07921__727 VPWR VGND net727 sg13g2_tiehi
XFILLER_7_996 VPWR VGND sg13g2_decap_8
XFILLER_43_4 VPWR VGND sg13g2_decap_4
XFILLER_97_712 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_181_clk_regs clknet_5_3__leaf_clk_regs clknet_leaf_181_clk_regs VPWR
+ VGND sg13g2_buf_8
Xhold1608 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[22\]
+ VPWR VGND net3435 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_110_clk_regs clknet_5_25__leaf_clk_regs clknet_leaf_110_clk_regs VPWR
+ VGND sg13g2_buf_8
X_07750_ net3256 net3270 net989 _01235_ VPWR VGND sg13g2_mux2_1
X_08234__443 VPWR VGND net443 sg13g2_tiehi
Xhold1619 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[19\]
+ VPWR VGND net3446 sg13g2_dlygate4sd3_1
X_04962_ _01693_ VPWR _01694_ VGND i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[1\]
+ _01688_ sg13g2_o21ai_1
X_08597__1379 VPWR VGND net1799 sg13g2_tiehi
X_06701_ VGND VPWR _02733_ _02736_ _02737_ net1181 sg13g2_a21oi_1
X_08771__1217 VPWR VGND net1637 sg13g2_tiehi
Xclkbuf_4_9_0_clk_regs clknet_0_clk_regs clknet_4_9_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_93_984 VPWR VGND sg13g2_decap_8
X_08089__605 VPWR VGND net605 sg13g2_tiehi
X_07681_ net2420 net3238 net1000 _01183_ VPWR VGND sg13g2_mux2_1
X_04893_ net1223 _01613_ _01616_ _01625_ VPWR VGND sg13g2_nor3_2
X_06632_ net1974 net1154 _02678_ VPWR VGND sg13g2_nor2_1
X_06563_ net3493 net1152 _02632_ VPWR VGND sg13g2_nor2_1
X_08302_ net376 VGND VPWR _00383_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[4\]
+ clknet_leaf_83_clk_regs sg13g2_dfrbpq_1
X_09282_ net57 VGND VPWR net2685 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[8\]
+ clknet_leaf_175_clk_regs sg13g2_dfrbpq_1
X_05514_ _02203_ VPWR i_exotiny._1611_\[18\] VGND net1074 _02205_ sg13g2_o21ai_1
X_08233_ net444 VGND VPWR net3128 i_exotiny._0028_\[0\] clknet_leaf_56_clk_regs sg13g2_dfrbpq_2
X_06494_ net2583 net3101 net1027 _00575_ VPWR VGND sg13g2_mux2_1
X_08241__436 VPWR VGND net436 sg13g2_tiehi
X_05445_ _02153_ VPWR net27 VGND i_exotiny._1660_ _01403_ sg13g2_o21ai_1
X_05376_ net1263 _01402_ _02076_ _02098_ VPWR VGND sg13g2_nor3_1
X_08164_ net514 VGND VPWR net2589 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[28\]
+ clknet_leaf_119_clk_regs sg13g2_dfrbpq_1
X_07115_ net1289 net1855 _00865_ VPWR VGND sg13g2_and2_1
X_08095_ net599 VGND VPWR net3418 i_exotiny._0013_\[0\] clknet_leaf_124_clk_regs sg13g2_dfrbpq_2
XFILLER_106_349 VPWR VGND sg13g2_decap_8
X_07046_ net2393 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[12\]
+ net1013 _00807_ VPWR VGND sg13g2_mux2_1
X_08419__266 VPWR VGND net266 sg13g2_tiehi
XFILLER_102_511 VPWR VGND sg13g2_decap_8
XFILLER_88_778 VPWR VGND sg13g2_fill_1
XFILLER_87_255 VPWR VGND sg13g2_fill_1
XFILLER_69_970 VPWR VGND sg13g2_fill_1
X_08997_ net1405 VGND VPWR net3566 i_exotiny._1160_\[18\] clknet_leaf_162_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_47_119 VPWR VGND sg13g2_fill_1
X_08747__1241 VPWR VGND net1661 sg13g2_tiehi
X_07948_ net708 VGND VPWR _00013_ i_exotiny._1623_ clknet_leaf_21_clk_regs sg13g2_dfrbpq_2
X_07879_ net2211 net2981 net978 _01346_ VPWR VGND sg13g2_mux2_1
X_08426__259 VPWR VGND net259 sg13g2_tiehi
XFILLER_34_43 VPWR VGND sg13g2_fill_2
XFILLER_8_738 VPWR VGND sg13g2_fill_2
XFILLER_11_288 VPWR VGND sg13g2_fill_1
X_08969__1013 VPWR VGND net1433 sg13g2_tiehi
XFILLER_50_75 VPWR VGND sg13g2_fill_1
XFILLER_4_911 VPWR VGND sg13g2_decap_8
XFILLER_98_509 VPWR VGND sg13g2_decap_8
XFILLER_4_988 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_105_382 VPWR VGND sg13g2_decap_8
Xfanout1200 net3242 net1200 VPWR VGND sg13g2_buf_8
Xfanout1222 net1223 net1222 VPWR VGND sg13g2_buf_8
Xfanout1211 net1212 net1211 VPWR VGND sg13g2_buf_8
Xfanout1255 net1257 net1255 VPWR VGND sg13g2_buf_8
Xfanout1233 i_exotiny._0315_\[2\] net1233 VPWR VGND sg13g2_buf_8
Xfanout1244 net3767 net1244 VPWR VGND sg13g2_buf_1
Xfanout1288 net1289 net1288 VPWR VGND sg13g2_buf_2
XFILLER_93_247 VPWR VGND sg13g2_fill_1
Xfanout1277 net1278 net1277 VPWR VGND sg13g2_buf_8
Xfanout1266 net1267 net1266 VPWR VGND sg13g2_buf_8
XFILLER_74_472 VPWR VGND sg13g2_decap_4
XFILLER_35_837 VPWR VGND sg13g2_fill_2
XFILLER_90_954 VPWR VGND sg13g2_decap_8
XFILLER_91_93 VPWR VGND sg13g2_fill_2
XFILLER_61_199 VPWR VGND sg13g2_fill_2
XFILLER_30_597 VPWR VGND sg13g2_fill_2
X_05230_ _01958_ _01649_ i_exotiny._0042_\[1\] _01641_ i_exotiny._0035_\[1\] VPWR
+ VGND sg13g2_a22oi_1
X_05161_ _01891_ _01650_ i_exotiny._0016_\[2\] _01636_ i_exotiny._0019_\[2\] VPWR
+ VGND sg13g2_a22oi_1
X_08825__1163 VPWR VGND net1583 sg13g2_tiehi
Xhold727 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[24\]
+ VPWR VGND net2554 sg13g2_dlygate4sd3_1
Xhold705 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[29\]
+ VPWR VGND net2532 sg13g2_dlygate4sd3_1
Xhold716 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[21\]
+ VPWR VGND net2543 sg13g2_dlygate4sd3_1
Xhold749 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[29\]
+ VPWR VGND net2576 sg13g2_dlygate4sd3_1
Xhold738 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[6\]
+ VPWR VGND net2565 sg13g2_dlygate4sd3_1
X_05092_ net1245 net1254 _01422_ _01823_ VPWR VGND sg13g2_nor3_1
X_08271__407 VPWR VGND net407 sg13g2_tiehi
X_08920_ net1482 VGND VPWR _00978_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[18\]
+ clknet_leaf_63_clk_regs sg13g2_dfrbpq_1
X_08988__994 VPWR VGND net1414 sg13g2_tiehi
X_08851_ net1555 VGND VPWR net2053 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[18\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
Xhold1405 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[28\]
+ VPWR VGND net3232 sg13g2_dlygate4sd3_1
Xhold1416 i_exotiny._0314_\[19\] VPWR VGND net3243 sg13g2_dlygate4sd3_1
X_07802_ net2869 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[20\]
+ net893 _01281_ VPWR VGND sg13g2_mux2_1
Xhold1449 _00817_ VPWR VGND net3276 sg13g2_dlygate4sd3_1
X_05994_ net2343 net2754 net1050 _00196_ VPWR VGND sg13g2_mux2_1
Xhold1438 _00198_ VPWR VGND net3265 sg13g2_dlygate4sd3_1
X_08782_ net1626 VGND VPWR _00840_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[13\]
+ clknet_leaf_170_clk_regs sg13g2_dfrbpq_1
Xhold1427 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[17\]
+ VPWR VGND net3254 sg13g2_dlygate4sd3_1
X_07733_ net3075 net881 _03199_ _03202_ VPWR VGND sg13g2_mux2_1
X_04945_ net1109 _01676_ _01677_ VPWR VGND sg13g2_and2_1
XFILLER_81_932 VPWR VGND sg13g2_fill_2
XFILLER_66_995 VPWR VGND sg13g2_fill_1
X_07664_ _03193_ net1138 net1165 _03194_ VPWR VGND sg13g2_a21o_2
X_04876_ _01606_ _01601_ _01466_ _01608_ VPWR VGND sg13g2_a21o_1
XFILLER_92_291 VPWR VGND sg13g2_decap_8
X_06615_ net1194 _02665_ _02666_ _00645_ VPWR VGND sg13g2_nor3_1
XFILLER_37_185 VPWR VGND sg13g2_fill_2
X_07595_ _03168_ net3607 _03166_ VPWR VGND sg13g2_xnor2_1
XFILLER_13_509 VPWR VGND sg13g2_fill_1
X_06546_ net2491 _02625_ net930 _00617_ VPWR VGND sg13g2_mux2_1
X_08995__987 VPWR VGND net1407 sg13g2_tiehi
X_06477_ net3297 net3351 net1024 _00558_ VPWR VGND sg13g2_mux2_1
X_09265_ net99 VGND VPWR net2537 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[23\]
+ clknet_leaf_130_clk_regs sg13g2_dfrbpq_1
X_09196_ net785 VGND VPWR _01251_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[18\]
+ clknet_leaf_79_clk_regs sg13g2_dfrbpq_1
X_05428_ _01384_ _02128_ _02134_ _02137_ VPWR VGND sg13g2_nor3_1
X_08216_ net461 VGND VPWR _00297_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[15\]
+ clknet_leaf_150_clk_regs sg13g2_dfrbpq_1
X_05359_ _02081_ _00020_ i_exotiny._2034_\[6\] VPWR VGND sg13g2_nand2_1
X_08147_ net531 VGND VPWR net2612 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[11\]
+ clknet_leaf_118_clk_regs sg13g2_dfrbpq_1
XFILLER_106_146 VPWR VGND sg13g2_decap_8
X_08078_ net616 VGND VPWR _00159_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[15\]
+ clknet_leaf_92_clk_regs sg13g2_dfrbpq_1
XFILLER_1_936 VPWR VGND sg13g2_decap_8
X_07029_ net3077 _02932_ net919 _00793_ VPWR VGND sg13g2_mux2_1
XFILLER_103_853 VPWR VGND sg13g2_decap_8
X_07994__135 VPWR VGND net135 sg13g2_tiehi
Xhold21 i_exotiny.i_wb_spi.state_r\[5\] VPWR VGND net1848 sg13g2_dlygate4sd3_1
Xhold10 i_exotiny.i_wb_spi.state_r\[13\] VPWR VGND net1837 sg13g2_dlygate4sd3_1
Xhold32 i_exotiny.i_wb_spi.state_r\[17\] VPWR VGND net1859 sg13g2_dlygate4sd3_1
XFILLER_49_918 VPWR VGND sg13g2_fill_2
XFILLER_102_385 VPWR VGND sg13g2_decap_8
Xhold54 _03179_ VPWR VGND net1881 sg13g2_dlygate4sd3_1
Xhold65 _01127_ VPWR VGND net1892 sg13g2_dlygate4sd3_1
Xhold43 i_exotiny.i_wdg_top.o_wb_dat\[11\] VPWR VGND net1870 sg13g2_dlygate4sd3_1
X_08217__460 VPWR VGND net460 sg13g2_tiehi
XFILLER_29_87 VPWR VGND sg13g2_fill_1
Xhold87 _03162_ VPWR VGND net1914 sg13g2_dlygate4sd3_1
Xhold1950 i_exotiny.i_wb_spi.dat_rx_r\[13\] VPWR VGND net3777 sg13g2_dlygate4sd3_1
Xhold76 i_exotiny._1924_\[3\] VPWR VGND net1903 sg13g2_dlygate4sd3_1
Xhold98 _00052_ VPWR VGND net1925 sg13g2_dlygate4sd3_1
Xhold1972 i_exotiny._1611_\[30\] VPWR VGND net3799 sg13g2_dlygate4sd3_1
Xhold1961 i_exotiny._6090_\[1\] VPWR VGND net3788 sg13g2_dlygate4sd3_1
Xhold1994 _02745_ VPWR VGND net3821 sg13g2_dlygate4sd3_1
Xhold1983 i_exotiny._0077_\[2\] VPWR VGND net3810 sg13g2_dlygate4sd3_1
XFILLER_72_943 VPWR VGND sg13g2_fill_2
XFILLER_45_53 VPWR VGND sg13g2_fill_2
XFILLER_71_486 VPWR VGND sg13g2_fill_2
XFILLER_71_453 VPWR VGND sg13g2_fill_2
X_07911__737 VPWR VGND net737 sg13g2_tiehi
X_08224__453 VPWR VGND net453 sg13g2_tiehi
XFILLER_8_535 VPWR VGND sg13g2_fill_2
X_08079__615 VPWR VGND net615 sg13g2_tiehi
XFILLER_98_306 VPWR VGND sg13g2_decap_8
XFILLER_4_785 VPWR VGND sg13g2_decap_8
Xfanout1030 net1031 net1030 VPWR VGND sg13g2_buf_8
XFILLER_6_1018 VPWR VGND sg13g2_decap_8
Xfanout1041 net1042 net1041 VPWR VGND sg13g2_buf_8
Xclkbuf_5_11__f_clk_regs clknet_4_5_0_clk_regs clknet_5_11__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
Xfanout1063 net1064 net1063 VPWR VGND sg13g2_buf_8
XFILLER_66_203 VPWR VGND sg13g2_fill_1
Xfanout1052 _02494_ net1052 VPWR VGND sg13g2_buf_8
XFILLER_0_980 VPWR VGND sg13g2_decap_8
Xfanout1074 net1075 net1074 VPWR VGND sg13g2_buf_8
Xfanout1096 net1101 net1096 VPWR VGND sg13g2_buf_8
XFILLER_54_409 VPWR VGND sg13g2_fill_2
X_08231__446 VPWR VGND net446 sg13g2_tiehi
Xfanout1085 _02990_ net1085 VPWR VGND sg13g2_buf_2
X_04730_ _01486_ net1230 net1231 VPWR VGND sg13g2_nand2_1
XFILLER_90_751 VPWR VGND sg13g2_fill_2
XFILLER_34_111 VPWR VGND sg13g2_fill_1
X_08086__608 VPWR VGND net608 sg13g2_tiehi
XFILLER_35_667 VPWR VGND sg13g2_fill_2
X_04661_ _01422_ _01420_ VPWR VGND net1247 sg13g2_nand2b_2
X_06400_ VGND VPWR net3778 _02180_ _02585_ net1225 sg13g2_a21oi_1
X_08409__276 VPWR VGND net276 sg13g2_tiehi
X_07380_ _03036_ _03025_ _03035_ net1210 i_exotiny._1160_\[8\] VPWR VGND sg13g2_a22oi_1
X_06331_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[29\]
+ net2730 net1034 _00468_ VPWR VGND sg13g2_mux2_1
X_06262_ net3231 net878 _02546_ _02550_ VPWR VGND sg13g2_mux2_1
X_09050_ net1352 VGND VPWR net1884 i_exotiny.i_rstctl.cnt\[0\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_2
X_08001_ net694 VGND VPWR _00082_ i_exotiny._0018_\[2\] clknet_leaf_69_clk_regs sg13g2_dfrbpq_2
X_05213_ VPWR VGND i_exotiny._0038_\[1\] _01940_ _01792_ i_exotiny._0014_\[1\] _01941_
+ _01760_ sg13g2_a221oi_1
X_06193_ net2230 i_exotiny._0033_\[1\] net945 _00348_ VPWR VGND sg13g2_mux2_1
Xhold502 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[18\]
+ VPWR VGND net2329 sg13g2_dlygate4sd3_1
Xhold524 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[18\]
+ VPWR VGND net2351 sg13g2_dlygate4sd3_1
Xhold513 _00974_ VPWR VGND net2340 sg13g2_dlygate4sd3_1
Xhold535 _00966_ VPWR VGND net2362 sg13g2_dlygate4sd3_1
X_05144_ _01874_ _01626_ i_exotiny._0014_\[2\] _01622_ i_exotiny._0023_\[2\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_104_628 VPWR VGND sg13g2_fill_2
Xhold579 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[22\]
+ VPWR VGND net2406 sg13g2_dlygate4sd3_1
Xhold546 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[21\]
+ VPWR VGND net2373 sg13g2_dlygate4sd3_1
Xhold557 _00439_ VPWR VGND net2384 sg13g2_dlygate4sd3_1
X_07978__119 VPWR VGND net119 sg13g2_tiehi
X_05075_ _01807_ _01788_ i_exotiny._0039_\[3\] _01769_ i_exotiny._0022_\[3\] VPWR
+ VGND sg13g2_a22oi_1
Xhold568 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[19\]
+ VPWR VGND net2395 sg13g2_dlygate4sd3_1
X_08903_ net1499 VGND VPWR net2890 i_exotiny._0040_\[1\] clknet_leaf_112_clk_regs
+ sg13g2_dfrbpq_2
X_09047__1151 VPWR VGND net1571 sg13g2_tiehi
XFILLER_100_812 VPWR VGND sg13g2_decap_8
XFILLER_85_501 VPWR VGND sg13g2_fill_2
X_08416__269 VPWR VGND net269 sg13g2_tiehi
Xhold1224 _01262_ VPWR VGND net3051 sg13g2_dlygate4sd3_1
XFILLER_98_895 VPWR VGND sg13g2_decap_8
XFILLER_97_394 VPWR VGND sg13g2_decap_8
Xhold1202 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[5\]
+ VPWR VGND net3029 sg13g2_dlygate4sd3_1
X_08834_ net1574 VGND VPWR net2205 i_exotiny._0036_\[1\] clknet_leaf_181_clk_regs
+ sg13g2_dfrbpq_2
Xhold1213 _00832_ VPWR VGND net3040 sg13g2_dlygate4sd3_1
X_08765_ net1643 VGND VPWR net3305 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[28\]
+ clknet_leaf_80_clk_regs sg13g2_dfrbpq_1
Xhold1257 _00962_ VPWR VGND net3084 sg13g2_dlygate4sd3_1
XFILLER_57_258 VPWR VGND sg13g2_decap_8
Xhold1246 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[6\]
+ VPWR VGND net3073 sg13g2_dlygate4sd3_1
Xhold1235 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[10\]
+ VPWR VGND net3062 sg13g2_dlygate4sd3_1
XFILLER_100_889 VPWR VGND sg13g2_decap_8
X_07716_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[17\]
+ net2579 net994 _01212_ VPWR VGND sg13g2_mux2_1
Xhold1268 _00588_ VPWR VGND net3095 sg13g2_dlygate4sd3_1
Xhold1279 _01135_ VPWR VGND net3106 sg13g2_dlygate4sd3_1
XFILLER_38_450 VPWR VGND sg13g2_fill_1
X_05977_ net2758 net3410 net1051 _00179_ VPWR VGND sg13g2_mux2_1
XFILLER_65_280 VPWR VGND sg13g2_fill_2
X_08696_ net1712 VGND VPWR net2926 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[23\]
+ clknet_leaf_105_clk_regs sg13g2_dfrbpq_1
X_04928_ _01660_ _01654_ i_exotiny._0020_\[3\] _01653_ i_exotiny._0038_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_04859_ VGND VPWR net1072 _01592_ i_exotiny._1902_\[5\] _01593_ sg13g2_a21oi_1
X_07647_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[20\]
+ net2236 net899 _01155_ VPWR VGND sg13g2_mux2_1
X_07578_ VGND VPWR i_exotiny.i_wdg_top.clk_div_inst.cnt\[2\] _03154_ _03157_ net1885
+ sg13g2_a21oi_1
XFILLER_13_328 VPWR VGND sg13g2_fill_2
X_06529_ net2184 net2437 net929 _00604_ VPWR VGND sg13g2_mux2_1
X_08697__1291 VPWR VGND net1711 sg13g2_tiehi
XFILLER_31_33 VPWR VGND sg13g2_decap_8
X_09248_ net559 VGND VPWR _01303_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[6\]
+ clknet_leaf_123_clk_regs sg13g2_dfrbpq_1
X_09179_ net802 VGND VPWR net2601 i_exotiny._0026_\[1\] clknet_leaf_80_clk_regs sg13g2_dfrbpq_2
X_08592__1384 VPWR VGND net1804 sg13g2_tiehi
Xoutput22 net22 uio_oe[4] VPWR VGND sg13g2_buf_1
Xoutput33 net33 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_733 VPWR VGND sg13g2_decap_8
XFILLER_103_661 VPWR VGND sg13g2_fill_1
XFILLER_102_182 VPWR VGND sg13g2_decap_8
XFILLER_76_556 VPWR VGND sg13g2_fill_1
Xhold1780 i_exotiny.i_wdg_top.clk_div_inst.cnt\[9\] VPWR VGND net3607 sg13g2_dlygate4sd3_1
XFILLER_63_217 VPWR VGND sg13g2_fill_2
Xhold1791 i_exotiny._2025_\[4\] VPWR VGND net3618 sg13g2_dlygate4sd3_1
XFILLER_72_51 VPWR VGND sg13g2_fill_2
XFILLER_44_486 VPWR VGND sg13g2_fill_2
XFILLER_12_372 VPWR VGND sg13g2_fill_1
XFILLER_8_321 VPWR VGND sg13g2_fill_2
XFILLER_40_692 VPWR VGND sg13g2_fill_2
XFILLER_4_582 VPWR VGND sg13g2_fill_1
X_08985__997 VPWR VGND net1417 sg13g2_tiehi
XFILLER_79_383 VPWR VGND sg13g2_fill_1
X_05900_ net2128 net2552 net972 _00117_ VPWR VGND sg13g2_mux2_1
X_06880_ VGND VPWR net1094 _02886_ _00689_ _02887_ sg13g2_a21oi_1
Xclkbuf_leaf_17_clk_regs clknet_5_6__leaf_clk_regs clknet_leaf_17_clk_regs VPWR VGND
+ sg13g2_buf_8
X_05831_ net2732 net2287 net1054 _00103_ VPWR VGND sg13g2_mux2_1
XFILLER_11_2 VPWR VGND sg13g2_fill_1
XFILLER_95_898 VPWR VGND sg13g2_decap_8
X_05762_ _02392_ VPWR _00066_ VGND net1143 _02391_ sg13g2_o21ai_1
X_08550_ net106 VGND VPWR _00624_ i_exotiny._0077_\[1\] clknet_leaf_160_clk_regs sg13g2_dfrbpq_1
X_08481_ net199 VGND VPWR _00555_ i_exotiny._0041_\[1\] clknet_leaf_70_clk_regs sg13g2_dfrbpq_2
X_05693_ net2528 net1064 _02341_ VPWR VGND sg13g2_nor2_1
X_07501_ i_exotiny._0315_\[18\] net3547 net905 _01084_ VPWR VGND sg13g2_mux2_1
X_04713_ _01461_ _01464_ _01466_ _01470_ _01471_ VPWR VGND sg13g2_nor4_1
XFILLER_74_1028 VPWR VGND sg13g2_fill_1
X_04644_ _01406_ net2997 VPWR VGND sg13g2_inv_2
X_07432_ net3387 net1214 _03076_ VPWR VGND sg13g2_and2_1
XFILLER_35_486 VPWR VGND sg13g2_fill_2
X_09102_ net1300 VGND VPWR _01157_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[22\]
+ clknet_leaf_144_clk_regs sg13g2_dfrbpq_1
X_07363_ _03023_ _03004_ _02629_ net1079 net3712 VPWR VGND sg13g2_a22oi_1
X_07294_ net2846 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[23\]
+ net911 _01011_ VPWR VGND sg13g2_mux2_1
X_06314_ net2325 net2426 net1036 _00451_ VPWR VGND sg13g2_mux2_1
X_08207__470 VPWR VGND net470 sg13g2_tiehi
X_06245_ net2939 net2914 net1039 _00394_ VPWR VGND sg13g2_mux2_1
XFILLER_11_1023 VPWR VGND sg13g2_decap_4
X_09033_ net1369 VGND VPWR _01091_ i_exotiny._0315_\[21\] clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
X_06176_ net2554 net2768 net953 _00338_ VPWR VGND sg13g2_mux2_1
Xhold310 _00382_ VPWR VGND net2137 sg13g2_dlygate4sd3_1
XFILLER_105_937 VPWR VGND sg13g2_decap_8
Xhold343 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[17\]
+ VPWR VGND net2170 sg13g2_dlygate4sd3_1
Xhold321 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[13\]
+ VPWR VGND net2148 sg13g2_dlygate4sd3_1
Xhold332 _00844_ VPWR VGND net2159 sg13g2_dlygate4sd3_1
X_05127_ _01857_ _01792_ i_exotiny._0038_\[2\] _01774_ i_exotiny._0018_\[2\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_104_425 VPWR VGND sg13g2_decap_8
Xhold354 _00397_ VPWR VGND net2181 sg13g2_dlygate4sd3_1
Xhold376 _00995_ VPWR VGND net2203 sg13g2_dlygate4sd3_1
Xhold387 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[7\]
+ VPWR VGND net2214 sg13g2_dlygate4sd3_1
Xhold365 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[24\]
+ VPWR VGND net2192 sg13g2_dlygate4sd3_1
Xhold398 _00601_ VPWR VGND net2225 sg13g2_dlygate4sd3_1
X_05058_ i_exotiny._0079_\[2\] i_exotiny._0079_\[3\] net1235 _01790_ VGND VPWR _01756_
+ sg13g2_nor4_2
X_08817_ net1591 VGND VPWR _00875_ i_exotiny.i_wb_spi.state_r\[16\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
Xhold1010 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[20\]
+ VPWR VGND net2837 sg13g2_dlygate4sd3_1
Xfanout889 net890 net889 VPWR VGND sg13g2_buf_8
Xfanout878 net879 net878 VPWR VGND sg13g2_buf_8
Xhold1032 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[11\]
+ VPWR VGND net2859 sg13g2_dlygate4sd3_1
Xhold1021 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[11\]
+ VPWR VGND net2848 sg13g2_dlygate4sd3_1
Xhold1076 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[15\]
+ VPWR VGND net2903 sg13g2_dlygate4sd3_1
Xhold1065 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[19\]
+ VPWR VGND net2892 sg13g2_dlygate4sd3_1
Xhold1054 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[9\]
+ VPWR VGND net2881 sg13g2_dlygate4sd3_1
Xhold1043 _01281_ VPWR VGND net2870 sg13g2_dlygate4sd3_1
X_08214__463 VPWR VGND net463 sg13g2_tiehi
X_08748_ net1660 VGND VPWR _00806_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[11\]
+ clknet_leaf_81_clk_regs sg13g2_dfrbpq_1
Xhold1087 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[15\]
+ VPWR VGND net2914 sg13g2_dlygate4sd3_1
Xhold1098 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[27\]
+ VPWR VGND net2925 sg13g2_dlygate4sd3_1
X_08069__625 VPWR VGND net625 sg13g2_tiehi
X_08679_ net1729 VGND VPWR _00737_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[6\]
+ clknet_leaf_103_clk_regs sg13g2_dfrbpq_1
XFILLER_54_773 VPWR VGND sg13g2_fill_2
XFILLER_54_762 VPWR VGND sg13g2_fill_1
X_09097__885 VPWR VGND net1305 sg13g2_tiehi
X_08784__1204 VPWR VGND net1624 sg13g2_tiehi
XFILLER_9_129 VPWR VGND sg13g2_fill_2
XFILLER_42_54 VPWR VGND sg13g2_decap_8
XFILLER_42_87 VPWR VGND sg13g2_fill_2
XFILLER_10_887 VPWR VGND sg13g2_fill_2
XFILLER_6_836 VPWR VGND sg13g2_decap_8
X_08221__456 VPWR VGND net456 sg13g2_tiehi
X_08076__618 VPWR VGND net618 sg13g2_tiehi
Xclkbuf_4_11_0_clk_regs clknet_0_clk_regs clknet_4_11_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_97_1028 VPWR VGND sg13g2_fill_1
XFILLER_97_1017 VPWR VGND sg13g2_decap_8
XFILLER_83_61 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_135_clk_regs clknet_5_21__leaf_clk_regs clknet_leaf_135_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_32_423 VPWR VGND sg13g2_fill_2
X_08406__279 VPWR VGND net279 sg13g2_tiehi
XFILLER_60_798 VPWR VGND sg13g2_fill_1
X_06030_ _02477_ _02509_ _02510_ VPWR VGND sg13g2_nor2_2
XFILLER_99_423 VPWR VGND sg13g2_decap_8
XFILLER_87_607 VPWR VGND sg13g2_fill_2
X_07981_ net122 VGND VPWR net3388 i_exotiny._0369_\[19\] clknet_leaf_14_clk_regs sg13g2_dfrbpq_2
X_06932_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[12\]
+ net3380 net926 _00711_ VPWR VGND sg13g2_mux2_1
XFILLER_41_1027 VPWR VGND sg13g2_fill_2
XFILLER_94_150 VPWR VGND sg13g2_fill_1
XFILLER_55_526 VPWR VGND sg13g2_fill_2
X_06863_ net3584 net1188 _02873_ VPWR VGND sg13g2_nor2_1
X_05814_ net2598 net2802 net1057 _00086_ VPWR VGND sg13g2_mux2_1
X_06794_ VGND VPWR net1098 _02814_ _00675_ _02815_ sg13g2_a21oi_1
X_08602_ net1794 VGND VPWR _00674_ i_exotiny._1615_\[2\] clknet_leaf_23_clk_regs sg13g2_dfrbpq_2
X_05745_ i_exotiny.i_wb_spi.cnt_hbit_r\[5\] net1930 _02368_ _02381_ VPWR VGND sg13g2_nor3_1
X_08533_ net147 VGND VPWR net2624 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[21\]
+ clknet_leaf_183_clk_regs sg13g2_dfrbpq_1
X_08905__1077 VPWR VGND net1497 sg13g2_tiehi
XFILLER_23_412 VPWR VGND sg13g2_fill_1
X_05676_ net1121 net1947 _02328_ VPWR VGND sg13g2_nor2b_1
X_08464_ net216 VGND VPWR net2738 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[16\]
+ clknet_leaf_64_clk_regs sg13g2_dfrbpq_1
XFILLER_50_220 VPWR VGND sg13g2_fill_2
XFILLER_35_294 VPWR VGND sg13g2_fill_1
X_04627_ VPWR _01389_ net3586 VGND sg13g2_inv_1
X_08395_ net535 VGND VPWR i_exotiny._1902_\[1\] i_exotiny.i_wb_spi.cnt_presc_r\[1\]
+ clknet_leaf_32_clk_regs sg13g2_dfrbpq_1
XFILLER_50_264 VPWR VGND sg13g2_fill_1
X_07415_ net1083 net3526 _03063_ _01048_ VPWR VGND sg13g2_a21o_1
X_07346_ _02992_ VPWR _03009_ VGND _02999_ _03004_ sg13g2_o21ai_1
X_07277_ net3168 net3210 net912 _00994_ VPWR VGND sg13g2_mux2_1
X_09016_ net1386 VGND VPWR _01074_ i_exotiny._0315_\[4\] clknet_leaf_9_clk_regs sg13g2_dfrbpq_2
X_06228_ _02525_ _02532_ _02546_ VPWR VGND sg13g2_nor2_2
XFILLER_105_734 VPWR VGND sg13g2_decap_8
XFILLER_104_222 VPWR VGND sg13g2_decap_8
X_06159_ net3102 net2739 net950 _00321_ VPWR VGND sg13g2_mux2_1
Xhold151 i_exotiny._1924_\[2\] VPWR VGND net1978 sg13g2_dlygate4sd3_1
Xhold140 i_exotiny.i_wb_spi.dat_rx_r\[5\] VPWR VGND net1967 sg13g2_dlygate4sd3_1
Xhold162 i_exotiny._1160_\[4\] VPWR VGND net1989 sg13g2_dlygate4sd3_1
Xhold173 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[23\]
+ VPWR VGND net2000 sg13g2_dlygate4sd3_1
Xhold195 i_exotiny._1160_\[8\] VPWR VGND net2022 sg13g2_dlygate4sd3_1
Xhold184 _01050_ VPWR VGND net2011 sg13g2_dlygate4sd3_1
XFILLER_104_299 VPWR VGND sg13g2_decap_8
XFILLER_101_962 VPWR VGND sg13g2_decap_8
XFILLER_58_353 VPWR VGND sg13g2_fill_2
XFILLER_100_472 VPWR VGND sg13g2_decap_8
XFILLER_37_43 VPWR VGND sg13g2_decap_4
XFILLER_37_65 VPWR VGND sg13g2_decap_4
XFILLER_73_345 VPWR VGND sg13g2_fill_1
XFILLER_6_600 VPWR VGND sg13g2_fill_2
XFILLER_97_905 VPWR VGND sg13g2_decap_8
XFILLER_69_618 VPWR VGND sg13g2_fill_1
XFILLER_96_437 VPWR VGND sg13g2_decap_8
XFILLER_78_83 VPWR VGND sg13g2_fill_1
XFILLER_2_894 VPWR VGND sg13g2_decap_8
XFILLER_37_504 VPWR VGND sg13g2_fill_1
XFILLER_64_378 VPWR VGND sg13g2_fill_1
XFILLER_60_540 VPWR VGND sg13g2_fill_2
X_05530_ _02215_ VPWR i_exotiny._1611_\[23\] VGND net1075 _02217_ sg13g2_o21ai_1
XFILLER_60_584 VPWR VGND sg13g2_fill_2
X_05461_ _02167_ VPWR net30 VGND net1264 _01404_ sg13g2_o21ai_1
X_05392_ net1112 _02109_ i_exotiny._2043_\[1\] VPWR VGND sg13g2_nor2_1
X_07200_ net1935 net1091 _02962_ VPWR VGND sg13g2_nor2_1
X_08180_ net497 VGND VPWR _00261_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[11\]
+ clknet_leaf_109_clk_regs sg13g2_dfrbpq_1
XFILLER_32_286 VPWR VGND sg13g2_fill_2
X_07131_ net1287 net1856 _00881_ VPWR VGND sg13g2_and2_1
XFILLER_64_0 VPWR VGND sg13g2_fill_1
X_07062_ i_exotiny._0017_\[0\] net888 _02934_ _02936_ VPWR VGND sg13g2_mux2_1
X_08204__473 VPWR VGND net473 sg13g2_tiehi
X_06013_ VGND VPWR net1980 net1106 _00209_ _02500_ sg13g2_a21oi_1
Xclkbuf_leaf_32_clk_regs clknet_5_8__leaf_clk_regs clknet_leaf_32_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08059__635 VPWR VGND net635 sg13g2_tiehi
X_09087__895 VPWR VGND net1315 sg13g2_tiehi
XFILLER_102_759 VPWR VGND sg13g2_decap_8
XFILLER_101_247 VPWR VGND sg13g2_decap_8
XFILLER_99_297 VPWR VGND sg13g2_decap_8
X_07964_ net1175 VGND VPWR net3797 i_exotiny.i_wdg_top.o_wb_dat\[5\] clknet_leaf_36_clk_regs
+ sg13g2_dfrbpq_1
X_06915_ _02914_ net2570 _02912_ VPWR VGND sg13g2_nand2_1
X_07895_ net3066 _03232_ net981 _01359_ VPWR VGND sg13g2_mux2_1
X_08586__740 VPWR VGND net740 sg13g2_tiehi
X_06846_ net1170 VPWR _02859_ VGND i_exotiny.i_wb_spi.dat_rx_r\[24\] net1186 sg13g2_o21ai_1
X_06777_ VGND VPWR _01415_ net1192 _02801_ net1169 sg13g2_a21oi_1
X_08211__466 VPWR VGND net466 sg13g2_tiehi
XFILLER_36_581 VPWR VGND sg13g2_fill_2
X_05728_ _02366_ net2033 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set[0]
+ _00058_ VPWR VGND sg13g2_a21o_1
X_08516_ net164 VGND VPWR net2836 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[4\]
+ clknet_leaf_176_clk_regs sg13g2_dfrbpq_1
X_08066__628 VPWR VGND net628 sg13g2_tiehi
X_08447_ net233 VGND VPWR _00521_ i_exotiny.i_wb_regs.spi_size_o\[1\] clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_2
X_05659_ net2004 net1063 _02315_ VPWR VGND sg13g2_nor2_1
X_09094__888 VPWR VGND net1308 sg13g2_tiehi
XFILLER_104_1021 VPWR VGND sg13g2_decap_8
X_08378_ net300 VGND VPWR net1977 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[16\]
+ clknet_leaf_137_clk_regs sg13g2_dfrbpq_1
XFILLER_20_982 VPWR VGND sg13g2_fill_1
X_07329_ _02993_ net1214 _02992_ VPWR VGND sg13g2_nand2_1
XFILLER_87_1027 VPWR VGND sg13g2_fill_2
XFILLER_105_564 VPWR VGND sg13g2_decap_8
X_08435__250 VPWR VGND net250 sg13g2_tiehi
XFILLER_87_971 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_64_41 VPWR VGND sg13g2_fill_1
X_08561__82 VPWR VGND net82 sg13g2_tiehi
XFILLER_11_960 VPWR VGND sg13g2_decap_8
X_08861__1125 VPWR VGND net1545 sg13g2_tiehi
XFILLER_7_975 VPWR VGND sg13g2_decap_8
Xhold909 i_exotiny._1611_\[29\] VPWR VGND net2736 sg13g2_dlygate4sd3_1
XFILLER_9_1027 VPWR VGND sg13g2_fill_2
XFILLER_9_1016 VPWR VGND sg13g2_decap_8
X_09305__933 VPWR VGND net1353 sg13g2_tiehi
XFILLER_97_757 VPWR VGND sg13g2_fill_1
Xhold1609 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[4\]
+ VPWR VGND net3436 sg13g2_dlygate4sd3_1
XFILLER_49_150 VPWR VGND sg13g2_fill_1
X_04961_ _01693_ _01363_ _01692_ VPWR VGND sg13g2_nand2_1
X_06700_ VGND VPWR i_exotiny._0369_\[1\] net1187 _02736_ net1219 sg13g2_a21oi_1
Xclkbuf_leaf_150_clk_regs clknet_5_16__leaf_clk_regs clknet_leaf_150_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_93_963 VPWR VGND sg13g2_decap_8
X_04892_ net1256 _01613_ _01623_ _01624_ VPWR VGND sg13g2_nor3_2
X_07680_ net2960 net3196 net998 _01182_ VPWR VGND sg13g2_mux2_1
X_06631_ i_exotiny._0314_\[23\] net1161 _02677_ VPWR VGND sg13g2_nor2_1
XFILLER_25_518 VPWR VGND sg13g2_fill_1
X_06562_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[0\].i_hadd.a_i
+ net1160 _02631_ VPWR VGND sg13g2_nor2_1
X_08301_ net377 VGND VPWR net2137 i_exotiny._0031_\[3\] clknet_leaf_73_clk_regs sg13g2_dfrbpq_2
X_09281_ net59 VGND VPWR net3141 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[7\]
+ clknet_leaf_171_clk_regs sg13g2_dfrbpq_1
X_05513_ VGND VPWR i_exotiny._0314_\[10\] net1276 _02205_ _02204_ sg13g2_a21oi_1
X_06493_ net2228 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[20\]
+ net1026 _00574_ VPWR VGND sg13g2_mux2_1
X_08232_ net445 VGND VPWR _00313_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[31\]
+ clknet_leaf_150_clk_regs sg13g2_dfrbpq_1
X_05444_ _02153_ _02151_ _02152_ VPWR VGND sg13g2_nand2b_1
X_05375_ net1263 _01402_ _02097_ VPWR VGND sg13g2_nor2_1
X_08163_ net515 VGND VPWR _00244_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[27\]
+ clknet_leaf_119_clk_regs sg13g2_dfrbpq_1
X_07114_ net1288 net1848 _00864_ VPWR VGND sg13g2_and2_1
X_08094_ net600 VGND VPWR net2506 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[31\]
+ clknet_leaf_85_clk_regs sg13g2_dfrbpq_1
XFILLER_106_328 VPWR VGND sg13g2_decap_8
X_07045_ net3199 net3449 net1016 _00806_ VPWR VGND sg13g2_mux2_1
X_09280__61 VPWR VGND net61 sg13g2_tiehi
XFILLER_0_606 VPWR VGND sg13g2_decap_4
XFILLER_0_628 VPWR VGND sg13g2_decap_4
XFILLER_102_534 VPWR VGND sg13g2_decap_8
X_08996_ net1406 VGND VPWR _01054_ i_exotiny._1160_\[17\] clknet_leaf_160_clk_regs
+ sg13g2_dfrbpq_1
X_07947_ net94 VGND VPWR _00012_ i_exotiny._1725_ clknet_leaf_22_clk_regs sg13g2_dfrbpq_2
XFILLER_28_301 VPWR VGND sg13g2_fill_1
XFILLER_55_142 VPWR VGND sg13g2_fill_1
X_07878_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[16\]
+ net2327 net979 _01345_ VPWR VGND sg13g2_mux2_1
XFILLER_28_356 VPWR VGND sg13g2_fill_1
XFILLER_84_996 VPWR VGND sg13g2_decap_8
XFILLER_83_484 VPWR VGND sg13g2_fill_2
XFILLER_83_473 VPWR VGND sg13g2_fill_1
X_06829_ net1132 _02843_ _02844_ _02845_ VPWR VGND sg13g2_nor3_1
X_08642__1335 VPWR VGND net1755 sg13g2_tiehi
XFILLER_34_66 VPWR VGND sg13g2_fill_2
XFILLER_4_967 VPWR VGND sg13g2_decap_8
XFILLER_106_895 VPWR VGND sg13g2_decap_8
XFILLER_105_361 VPWR VGND sg13g2_decap_8
XFILLER_78_234 VPWR VGND sg13g2_fill_1
Xfanout1201 _01434_ net1201 VPWR VGND sg13g2_buf_8
Xfanout1212 _01504_ net1212 VPWR VGND sg13g2_buf_8
Xfanout1223 _01394_ net1223 VPWR VGND sg13g2_buf_8
Xclkbuf_5_10__f_clk_regs clknet_4_5_0_clk_regs clknet_5_10__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08900__1082 VPWR VGND net1502 sg13g2_tiehi
Xfanout1234 net3688 net1234 VPWR VGND sg13g2_buf_8
Xfanout1256 net1257 net1256 VPWR VGND sg13g2_buf_8
Xfanout1245 i_exotiny._0542_ net1245 VPWR VGND sg13g2_buf_8
Xfanout1289 net1290 net1289 VPWR VGND sg13g2_buf_1
Xfanout1278 net1280 net1278 VPWR VGND sg13g2_buf_8
Xfanout1267 net3694 net1267 VPWR VGND sg13g2_buf_8
XFILLER_90_933 VPWR VGND sg13g2_decap_8
XFILLER_28_890 VPWR VGND sg13g2_fill_2
X_08049__645 VPWR VGND net645 sg13g2_tiehi
X_05160_ _01890_ _01645_ i_exotiny._0025_\[2\] _01637_ i_exotiny._0024_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold728 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[27\]
+ VPWR VGND net2555 sg13g2_dlygate4sd3_1
Xhold706 _00583_ VPWR VGND net2533 sg13g2_dlygate4sd3_1
Xhold717 _00101_ VPWR VGND net2544 sg13g2_dlygate4sd3_1
XFILLER_7_794 VPWR VGND sg13g2_fill_1
Xhold739 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[18\]
+ VPWR VGND net2566 sg13g2_dlygate4sd3_1
X_08201__476 VPWR VGND net476 sg13g2_tiehi
X_05091_ VGND VPWR _01822_ _01821_ _01680_ sg13g2_or2_1
X_08850_ net1556 VGND VPWR _00908_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[17\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
X_09084__898 VPWR VGND net1318 sg13g2_tiehi
XFILLER_97_587 VPWR VGND sg13g2_fill_2
XFILLER_97_554 VPWR VGND sg13g2_fill_2
Xhold1406 _01020_ VPWR VGND net3233 sg13g2_dlygate4sd3_1
X_08056__638 VPWR VGND net638 sg13g2_tiehi
Xclkbuf_5_29__f_clk_regs clknet_4_14_0_clk_regs clknet_5_29__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07801_ net2251 net3108 net891 _01280_ VPWR VGND sg13g2_mux2_1
Xhold1428 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[20\]
+ VPWR VGND net3255 sg13g2_dlygate4sd3_1
Xhold1439 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[19\]
+ VPWR VGND net3266 sg13g2_dlygate4sd3_1
Xhold1417 _00643_ VPWR VGND net3244 sg13g2_dlygate4sd3_1
X_08781_ net1627 VGND VPWR _00839_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[12\]
+ clknet_leaf_168_clk_regs sg13g2_dfrbpq_1
X_08720__1268 VPWR VGND net1688 sg13g2_tiehi
X_05993_ net2395 net2337 net1051 _00195_ VPWR VGND sg13g2_mux2_1
X_07732_ _03201_ net2839 net994 _01227_ VPWR VGND sg13g2_mux2_1
X_04944_ VGND VPWR _01675_ _01676_ _01612_ i_exotiny._0314_\[3\] sg13g2_a21oi_2
XFILLER_93_782 VPWR VGND sg13g2_fill_1
XFILLER_81_911 VPWR VGND sg13g2_fill_2
X_07663_ _02492_ _02532_ _03193_ VPWR VGND sg13g2_nor2_2
X_04875_ VGND VPWR _01466_ _01607_ _01606_ _01601_ sg13g2_a21oi_2
X_06614_ net3489 net1157 _02666_ VPWR VGND sg13g2_nor2_1
X_07594_ _03166_ _03167_ _01123_ VPWR VGND sg13g2_nor2_1
X_08425__260 VPWR VGND net260 sg13g2_tiehi
X_06545_ i_exotiny._0043_\[3\] net872 _02620_ _02625_ VPWR VGND sg13g2_mux2_1
X_06476_ net2081 i_exotiny._0041_\[3\] net1023 _00557_ VPWR VGND sg13g2_mux2_1
X_09264_ net101 VGND VPWR net3253 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[22\]
+ clknet_leaf_127_clk_regs sg13g2_dfrbpq_1
X_09195_ net786 VGND VPWR _01250_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[17\]
+ clknet_leaf_78_clk_regs sg13g2_dfrbpq_1
X_05427_ _01384_ _02134_ _02136_ VPWR VGND sg13g2_nor2_2
X_08215_ net462 VGND VPWR net3451 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[14\]
+ clknet_leaf_151_clk_regs sg13g2_dfrbpq_1
X_08146_ net539 VGND VPWR _00227_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[10\]
+ clknet_leaf_155_clk_regs sg13g2_dfrbpq_1
X_05358_ _00020_ i_exotiny._2034_\[6\] _02080_ VPWR VGND sg13g2_nor2_1
XFILLER_106_125 VPWR VGND sg13g2_decap_8
XFILLER_105_7 VPWR VGND sg13g2_fill_2
X_08077_ net617 VGND VPWR _00158_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[14\]
+ clknet_leaf_86_clk_regs sg13g2_dfrbpq_1
X_05289_ _02015_ _01621_ i_exotiny._0043_\[0\] _01619_ i_exotiny._0034_\[0\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_1_915 VPWR VGND sg13g2_decap_8
X_07028_ i_exotiny._0032_\[2\] net877 _02928_ _02932_ VPWR VGND sg13g2_mux2_1
XFILLER_103_832 VPWR VGND sg13g2_decap_8
Xhold11 i_exotiny.i_wb_spi.state_r\[27\] VPWR VGND net1838 sg13g2_dlygate4sd3_1
XFILLER_102_364 VPWR VGND sg13g2_decap_8
Xhold22 i_exotiny.i_wb_spi.state_r\[12\] VPWR VGND net1849 sg13g2_dlygate4sd3_1
X_08432__253 VPWR VGND net253 sg13g2_tiehi
Xhold55 _01131_ VPWR VGND net1882 sg13g2_dlygate4sd3_1
Xhold33 _00876_ VPWR VGND net1860 sg13g2_dlygate4sd3_1
Xhold44 _00077_ VPWR VGND net1871 sg13g2_dlygate4sd3_1
X_08979_ net1423 VGND VPWR _01037_ i_exotiny._1160_\[0\] clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
Xhold88 _01121_ VPWR VGND net1915 sg13g2_dlygate4sd3_1
Xhold77 _00028_ VPWR VGND net1904 sg13g2_dlygate4sd3_1
Xhold99 i_exotiny._1924_\[22\] VPWR VGND net1926 sg13g2_dlygate4sd3_1
Xhold1962 i_exotiny._0327_\[0\] VPWR VGND net3789 sg13g2_dlygate4sd3_1
Xhold66 i_exotiny._1429_ VPWR VGND net1893 sg13g2_dlygate4sd3_1
Xhold1940 i_exotiny._0601_ VPWR VGND net3767 sg13g2_dlygate4sd3_1
Xhold1951 i_exotiny._0369_\[8\] VPWR VGND net3778 sg13g2_dlygate4sd3_1
Xhold1973 i_exotiny._0369_\[5\] VPWR VGND net3800 sg13g2_dlygate4sd3_1
Xhold1995 i_exotiny._0315_\[6\] VPWR VGND net3822 sg13g2_dlygate4sd3_1
Xhold1984 i_exotiny._1618_\[0\] VPWR VGND net3811 sg13g2_dlygate4sd3_1
XFILLER_45_87 VPWR VGND sg13g2_fill_2
XFILLER_45_98 VPWR VGND sg13g2_decap_4
XFILLER_12_510 VPWR VGND sg13g2_fill_1
XFILLER_101_93 VPWR VGND sg13g2_fill_1
XFILLER_12_543 VPWR VGND sg13g2_fill_1
X_08918__1064 VPWR VGND net1484 sg13g2_tiehi
XFILLER_6_15 VPWR VGND sg13g2_fill_1
XFILLER_106_692 VPWR VGND sg13g2_decap_8
Xfanout1031 net1032 net1031 VPWR VGND sg13g2_buf_8
Xfanout1020 net1022 net1020 VPWR VGND sg13g2_buf_8
XFILLER_94_535 VPWR VGND sg13g2_decap_8
Xfanout1042 _02547_ net1042 VPWR VGND sg13g2_buf_8
Xfanout1064 net1067 net1064 VPWR VGND sg13g2_buf_2
Xfanout1053 net1055 net1053 VPWR VGND sg13g2_buf_8
Xfanout1086 net1091 net1086 VPWR VGND sg13g2_buf_8
Xfanout1097 net1099 net1097 VPWR VGND sg13g2_buf_8
Xfanout1075 net1076 net1075 VPWR VGND sg13g2_buf_8
XFILLER_35_635 VPWR VGND sg13g2_decap_4
X_04660_ net1247 _01420_ _01421_ VPWR VGND sg13g2_nor2b_2
X_06330_ net3223 net2429 net1035 _00467_ VPWR VGND sg13g2_mux2_1
X_06261_ _02549_ net3164 net1039 _00408_ VPWR VGND sg13g2_mux2_1
X_08000_ net695 VGND VPWR net2816 i_exotiny._0018_\[1\] clknet_leaf_69_clk_regs sg13g2_dfrbpq_2
X_05212_ _01927_ _01939_ _01922_ _01940_ VPWR VGND sg13g2_nand3_1
X_06192_ net2146 i_exotiny._0033_\[0\] net948 _00347_ VPWR VGND sg13g2_mux2_1
Xhold525 _00126_ VPWR VGND net2352 sg13g2_dlygate4sd3_1
Xhold514 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[30\]
+ VPWR VGND net2341 sg13g2_dlygate4sd3_1
Xhold536 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[27\]
+ VPWR VGND net2363 sg13g2_dlygate4sd3_1
Xhold503 _00745_ VPWR VGND net2330 sg13g2_dlygate4sd3_1
X_05143_ _01873_ _01642_ i_exotiny._0015_\[2\] _01630_ i_exotiny._0041_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold547 _00400_ VPWR VGND net2374 sg13g2_dlygate4sd3_1
Xhold558 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[11\]
+ VPWR VGND net2385 sg13g2_dlygate4sd3_1
Xhold569 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[25\]
+ VPWR VGND net2396 sg13g2_dlygate4sd3_1
X_05074_ VPWR VGND i_exotiny._0028_\[3\] _01805_ _01781_ i_exotiny._0032_\[3\] _01806_
+ _01767_ sg13g2_a221oi_1
X_08902_ net1500 VGND VPWR _00960_ i_exotiny._0040_\[0\] clknet_leaf_113_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_106_38 VPWR VGND sg13g2_decap_8
XFILLER_98_874 VPWR VGND sg13g2_decap_8
XFILLER_97_373 VPWR VGND sg13g2_decap_8
Xhold1203 _00145_ VPWR VGND net3030 sg13g2_dlygate4sd3_1
X_08833_ net1575 VGND VPWR net2175 i_exotiny._0036_\[0\] clknet_leaf_183_clk_regs
+ sg13g2_dfrbpq_2
Xhold1214 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[19\]
+ VPWR VGND net3041 sg13g2_dlygate4sd3_1
Xhold1225 i_exotiny._0315_\[27\] VPWR VGND net3052 sg13g2_dlygate4sd3_1
XFILLER_100_868 VPWR VGND sg13g2_decap_8
X_08764_ net1644 VGND VPWR _00822_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[27\]
+ clknet_leaf_81_clk_regs sg13g2_dfrbpq_1
X_05976_ i_exotiny._0013_\[2\] net2207 net1049 _00178_ VPWR VGND sg13g2_mux2_1
Xhold1258 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[28\]
+ VPWR VGND net3085 sg13g2_dlygate4sd3_1
Xhold1236 i_exotiny._0015_\[0\] VPWR VGND net3063 sg13g2_dlygate4sd3_1
Xhold1247 _00833_ VPWR VGND net3074 sg13g2_dlygate4sd3_1
XFILLER_38_440 VPWR VGND sg13g2_fill_1
X_09199__782 VPWR VGND net782 sg13g2_tiehi
Xhold1269 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[21\]
+ VPWR VGND net3096 sg13g2_dlygate4sd3_1
X_07715_ net2916 net2335 net993 _01211_ VPWR VGND sg13g2_mux2_1
X_04927_ _01639_ _01656_ _01633_ _01659_ VPWR VGND _01658_ sg13g2_nand4_1
XFILLER_66_793 VPWR VGND sg13g2_fill_1
X_08695_ net1713 VGND VPWR net2771 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[22\]
+ clknet_leaf_105_clk_regs sg13g2_dfrbpq_1
X_04858_ VGND VPWR net3561 _01570_ _01593_ net1072 sg13g2_a21oi_1
XFILLER_54_977 VPWR VGND sg13g2_fill_2
X_07646_ net2952 net3070 net896 _01154_ VPWR VGND sg13g2_mux2_1
XFILLER_25_156 VPWR VGND sg13g2_fill_1
X_07577_ VPWR _01117_ _03156_ VGND sg13g2_inv_1
X_04789_ _01539_ _01531_ _01535_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_104 VPWR VGND sg13g2_decap_4
XFILLER_41_638 VPWR VGND sg13g2_fill_2
XFILLER_41_649 VPWR VGND sg13g2_fill_2
X_06528_ net3054 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[21\]
+ net931 _00603_ VPWR VGND sg13g2_mux2_1
X_09247_ net560 VGND VPWR net3125 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[5\]
+ clknet_leaf_128_clk_regs sg13g2_dfrbpq_1
X_06459_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[28\]
+ net3151 net938 _00546_ VPWR VGND sg13g2_mux2_1
X_09178_ net803 VGND VPWR net3158 i_exotiny._0026_\[0\] clknet_leaf_78_clk_regs sg13g2_dfrbpq_2
X_08129_ net1177 VGND VPWR net2332 _00017_ clknet_leaf_36_clk_regs sg13g2_dfrbpq_2
Xoutput23 net23 uio_oe[5] VPWR VGND sg13g2_buf_1
Xoutput34 net34 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_0_244 VPWR VGND sg13g2_fill_2
XFILLER_103_673 VPWR VGND sg13g2_decap_4
X_08039__655 VPWR VGND net655 sg13g2_tiehi
X_08609__1367 VPWR VGND net1787 sg13g2_tiehi
XFILLER_1_789 VPWR VGND sg13g2_decap_8
XFILLER_56_53 VPWR VGND sg13g2_fill_2
Xhold1770 i_exotiny._1611_\[27\] VPWR VGND net3597 sg13g2_dlygate4sd3_1
Xhold1781 _03168_ VPWR VGND net3608 sg13g2_dlygate4sd3_1
Xhold1792 i_exotiny._1902_\[4\] VPWR VGND net3619 sg13g2_dlygate4sd3_1
XFILLER_71_262 VPWR VGND sg13g2_fill_2
XFILLER_13_863 VPWR VGND sg13g2_fill_1
X_08046__648 VPWR VGND net648 sg13g2_tiehi
XFILLER_82_9 VPWR VGND sg13g2_fill_2
XFILLER_67_1025 VPWR VGND sg13g2_decap_4
X_08092__602 VPWR VGND net602 sg13g2_tiehi
X_08415__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_95_877 VPWR VGND sg13g2_decap_8
X_05830_ net2666 net2504 net1054 _00102_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_57_clk_regs clknet_5_14__leaf_clk_regs clknet_leaf_57_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_67_579 VPWR VGND sg13g2_fill_1
XFILLER_48_771 VPWR VGND sg13g2_fill_2
X_05761_ _02392_ net1126 net3326 net1144 net3735 VPWR VGND sg13g2_a22oi_1
XFILLER_75_590 VPWR VGND sg13g2_fill_1
X_07500_ i_exotiny._0315_\[17\] net3545 net904 _01083_ VPWR VGND sg13g2_mux2_1
X_08480_ net200 VGND VPWR _00554_ i_exotiny._0041_\[0\] clknet_leaf_109_clk_regs sg13g2_dfrbpq_2
X_05692_ VGND VPWR i_exotiny._1616_\[3\] net1123 _02340_ _02339_ sg13g2_a21oi_1
X_04712_ i_exotiny._0571_ net1253 _01468_ _01470_ VPWR VGND sg13g2_nor3_2
XFILLER_62_284 VPWR VGND sg13g2_fill_1
X_04643_ VPWR _01405_ net12 VGND sg13g2_inv_1
XFILLER_23_638 VPWR VGND sg13g2_fill_1
X_07431_ net1081 net2020 _03075_ _01052_ VPWR VGND sg13g2_a21o_1
XFILLER_23_649 VPWR VGND sg13g2_fill_2
X_07362_ _03022_ _03009_ _03021_ net1208 net1989 VPWR VGND sg13g2_a22oi_1
X_09101_ net1301 VGND VPWR net2397 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[21\]
+ clknet_leaf_143_clk_regs sg13g2_dfrbpq_1
X_06313_ net2826 net3263 net1033 _00450_ VPWR VGND sg13g2_mux2_1
X_08422__263 VPWR VGND net263 sg13g2_tiehi
X_07293_ net2035 net3036 net909 _01010_ VPWR VGND sg13g2_mux2_1
X_06244_ net3285 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[14\]
+ net1038 _00393_ VPWR VGND sg13g2_mux2_1
XFILLER_11_1002 VPWR VGND sg13g2_decap_8
X_09032_ net1370 VGND VPWR net2842 i_exotiny._0315_\[20\] clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
Xhold300 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[17\]
+ VPWR VGND net2127 sg13g2_dlygate4sd3_1
Xhold311 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[4\]
+ VPWR VGND net2138 sg13g2_dlygate4sd3_1
X_06175_ net2238 net2591 net950 _00337_ VPWR VGND sg13g2_mux2_1
XFILLER_105_916 VPWR VGND sg13g2_decap_8
XFILLER_104_404 VPWR VGND sg13g2_decap_8
Xhold344 _00157_ VPWR VGND net2171 sg13g2_dlygate4sd3_1
Xhold333 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[30\]
+ VPWR VGND net2160 sg13g2_dlygate4sd3_1
Xhold322 _00259_ VPWR VGND net2149 sg13g2_dlygate4sd3_1
X_05126_ _01856_ _01788_ i_exotiny._0039_\[2\] _01758_ i_exotiny._0040_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold366 _00719_ VPWR VGND net2193 sg13g2_dlygate4sd3_1
Xhold377 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[5\]
+ VPWR VGND net2204 sg13g2_dlygate4sd3_1
Xhold355 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[4\]
+ VPWR VGND net2182 sg13g2_dlygate4sd3_1
Xhold399 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[25\]
+ VPWR VGND net2226 sg13g2_dlygate4sd3_1
Xhold388 _00083_ VPWR VGND net2215 sg13g2_dlygate4sd3_1
X_05057_ net1238 net1240 net1220 _01789_ VGND VPWR _01757_ sg13g2_nor4_2
Xhold1000 _00454_ VPWR VGND net2827 sg13g2_dlygate4sd3_1
Xhold1011 _01253_ VPWR VGND net2838 sg13g2_dlygate4sd3_1
X_08816_ net1592 VGND VPWR net1842 i_exotiny.i_wb_spi.state_r\[15\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
Xfanout879 net880 net879 VPWR VGND sg13g2_buf_8
Xhold1022 _00710_ VPWR VGND net2849 sg13g2_dlygate4sd3_1
Xhold1033 _01142_ VPWR VGND net2860 sg13g2_dlygate4sd3_1
Xhold1044 i_exotiny._0033_\[1\] VPWR VGND net2871 sg13g2_dlygate4sd3_1
Xhold1066 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[10\]
+ VPWR VGND net2893 sg13g2_dlygate4sd3_1
Xhold1055 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[11\]
+ VPWR VGND net2882 sg13g2_dlygate4sd3_1
X_05959_ net2234 net2812 net968 _00168_ VPWR VGND sg13g2_mux2_1
Xhold1077 _00123_ VPWR VGND net2904 sg13g2_dlygate4sd3_1
XFILLER_85_398 VPWR VGND sg13g2_fill_1
Xhold1088 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[26\]
+ VPWR VGND net2915 sg13g2_dlygate4sd3_1
X_08747_ net1661 VGND VPWR _00805_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[10\]
+ clknet_leaf_84_clk_regs sg13g2_dfrbpq_1
Xhold1099 _00754_ VPWR VGND net2926 sg13g2_dlygate4sd3_1
XFILLER_45_229 VPWR VGND sg13g2_fill_2
X_08678_ net1730 VGND VPWR _00736_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[5\]
+ clknet_leaf_112_clk_regs sg13g2_dfrbpq_1
X_07629_ i_exotiny._0024_\[2\] net2462 net897 _01137_ VPWR VGND sg13g2_mux2_1
XFILLER_42_925 VPWR VGND sg13g2_decap_4
XFILLER_14_649 VPWR VGND sg13g2_fill_2
XFILLER_50_991 VPWR VGND sg13g2_fill_1
XFILLER_6_826 VPWR VGND sg13g2_fill_1
XFILLER_6_804 VPWR VGND sg13g2_fill_2
XFILLER_96_619 VPWR VGND sg13g2_fill_1
XFILLER_104_993 VPWR VGND sg13g2_decap_8
XFILLER_77_866 VPWR VGND sg13g2_fill_2
XFILLER_49_535 VPWR VGND sg13g2_fill_2
XFILLER_92_803 VPWR VGND sg13g2_fill_2
XFILLER_91_302 VPWR VGND sg13g2_fill_2
XFILLER_91_368 VPWR VGND sg13g2_fill_1
XFILLER_60_755 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_175_clk_regs clknet_5_4__leaf_clk_regs clknet_leaf_175_clk_regs VPWR
+ VGND sg13g2_buf_8
Xclkbuf_leaf_104_clk_regs clknet_5_22__leaf_clk_regs clknet_leaf_104_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_8_152 VPWR VGND sg13g2_fill_1
X_08991__991 VPWR VGND net1411 sg13g2_tiehi
X_09189__792 VPWR VGND net792 sg13g2_tiehi
XFILLER_9_697 VPWR VGND sg13g2_fill_1
X_08376__302 VPWR VGND net302 sg13g2_tiehi
XFILLER_99_402 VPWR VGND sg13g2_decap_8
X_08655__1322 VPWR VGND net1742 sg13g2_tiehi
XFILLER_99_479 VPWR VGND sg13g2_decap_8
X_07980_ net121 VGND VPWR net3458 i_exotiny._0369_\[18\] clknet_leaf_13_clk_regs sg13g2_dfrbpq_2
XFILLER_101_429 VPWR VGND sg13g2_decap_8
X_06931_ net2848 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[15\]
+ net927 _00710_ VPWR VGND sg13g2_mux2_1
X_08601_ net1795 VGND VPWR _00673_ i_exotiny._1615_\[1\] clknet_leaf_24_clk_regs sg13g2_dfrbpq_2
X_06862_ VGND VPWR net1095 _02871_ _00686_ _02872_ sg13g2_a21oi_1
XFILLER_83_836 VPWR VGND sg13g2_fill_2
X_05813_ net2321 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[5\]
+ net1056 _00085_ VPWR VGND sg13g2_mux2_1
X_06793_ net3801 net1098 _02815_ VPWR VGND sg13g2_nor2_1
X_09196__785 VPWR VGND net785 sg13g2_tiehi
X_08877__1105 VPWR VGND net1525 sg13g2_tiehi
X_05744_ net1930 VPWR _02380_ VGND _01584_ _02379_ sg13g2_o21ai_1
X_08532_ net148 VGND VPWR _00606_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[20\]
+ clknet_leaf_176_clk_regs sg13g2_dfrbpq_1
X_08463_ net217 VGND VPWR _00537_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[15\]
+ clknet_leaf_159_clk_regs sg13g2_dfrbpq_1
X_05675_ net1957 net1062 _02327_ VPWR VGND sg13g2_nor2_1
X_07414_ net1083 _03061_ _03062_ _03063_ VPWR VGND sg13g2_nor3_1
X_08394_ net534 VGND VPWR i_exotiny._1902_\[0\] i_exotiny.i_wb_spi.cnt_presc_r\[0\]
+ clknet_leaf_32_clk_regs sg13g2_dfrbpq_2
X_04626_ net1268 _01388_ VPWR VGND sg13g2_inv_4
X_08029__665 VPWR VGND net665 sg13g2_tiehi
X_07345_ net2125 net1214 _03008_ VPWR VGND sg13g2_and2_1
X_07276_ net2840 net2654 net912 _00993_ VPWR VGND sg13g2_mux2_1
X_06227_ _02545_ net3208 net946 _00378_ VPWR VGND sg13g2_mux2_1
X_09015_ net1387 VGND VPWR _01073_ i_exotiny._0315_\[3\] clknet_leaf_9_clk_regs sg13g2_dfrbpq_2
XFILLER_105_713 VPWR VGND sg13g2_decap_8
XFILLER_104_201 VPWR VGND sg13g2_decap_8
X_06158_ net2166 net2557 net952 _00320_ VPWR VGND sg13g2_mux2_1
Xhold141 i_exotiny.i_wb_spi.dat_rx_r\[7\] VPWR VGND net1968 sg13g2_dlygate4sd3_1
Xhold130 i_exotiny._1924_\[20\] VPWR VGND net1957 sg13g2_dlygate4sd3_1
Xhold152 _00027_ VPWR VGND net1979 sg13g2_dlygate4sd3_1
Xhold185 i_exotiny._1614_\[1\] VPWR VGND net2012 sg13g2_dlygate4sd3_1
X_06089_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[15\]
+ net2073 net960 _00265_ VPWR VGND sg13g2_mux2_1
Xhold174 _00462_ VPWR VGND net2001 sg13g2_dlygate4sd3_1
X_05109_ VGND VPWR _01743_ _01838_ _01839_ _01702_ sg13g2_a21oi_1
Xhold163 _01041_ VPWR VGND net1990 sg13g2_dlygate4sd3_1
XFILLER_104_278 VPWR VGND sg13g2_decap_8
Xhold196 _01045_ VPWR VGND net2023 sg13g2_dlygate4sd3_1
XFILLER_101_941 VPWR VGND sg13g2_decap_8
XFILLER_100_451 VPWR VGND sg13g2_decap_8
X_08036__658 VPWR VGND net658 sg13g2_tiehi
XFILLER_18_207 VPWR VGND sg13g2_fill_2
XFILLER_37_11 VPWR VGND sg13g2_decap_4
XFILLER_74_869 VPWR VGND sg13g2_fill_2
XFILLER_15_925 VPWR VGND sg13g2_fill_1
XFILLER_26_262 VPWR VGND sg13g2_fill_2
XFILLER_42_700 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_2_clk_regs clknet_5_2__leaf_clk_regs clknet_leaf_2_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08733__1255 VPWR VGND net1675 sg13g2_tiehi
XFILLER_42_733 VPWR VGND sg13g2_fill_2
X_08082__612 VPWR VGND net612 sg13g2_tiehi
XFILLER_23_991 VPWR VGND sg13g2_fill_1
X_08405__280 VPWR VGND net280 sg13g2_tiehi
X_08955__1027 VPWR VGND net1447 sg13g2_tiehi
XFILLER_2_873 VPWR VGND sg13g2_decap_8
XFILLER_104_790 VPWR VGND sg13g2_decap_8
XFILLER_78_95 VPWR VGND sg13g2_fill_1
XFILLER_65_803 VPWR VGND sg13g2_fill_1
X_08412__273 VPWR VGND net273 sg13g2_tiehi
XFILLER_37_549 VPWR VGND sg13g2_decap_4
XFILLER_18_730 VPWR VGND sg13g2_decap_4
XFILLER_45_593 VPWR VGND sg13g2_fill_1
X_05460_ _02167_ _02165_ _02166_ VPWR VGND sg13g2_nand2b_1
X_05391_ _02109_ i_exotiny._2034_\[0\] i_exotiny._2034_\[1\] VPWR VGND sg13g2_xnor2_1
XFILLER_20_449 VPWR VGND sg13g2_fill_2
X_07130_ net1289 net1839 _00880_ VPWR VGND sg13g2_and2_1
X_07061_ net3047 net2555 net1015 _00822_ VPWR VGND sg13g2_mux2_1
X_08604__1372 VPWR VGND net1792 sg13g2_tiehi
X_06012_ _00016_ net1106 _02500_ VPWR VGND sg13g2_nor2_1
XFILLER_57_0 VPWR VGND sg13g2_fill_1
XFILLER_102_738 VPWR VGND sg13g2_decap_8
XFILLER_99_276 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_72_clk_regs clknet_5_27__leaf_clk_regs clknet_leaf_72_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08811__1177 VPWR VGND net1597 sg13g2_tiehi
XFILLER_101_226 VPWR VGND sg13g2_decap_8
X_07963_ net1175 VGND VPWR net3786 i_exotiny.i_wdg_top.o_wb_dat\[4\] clknet_leaf_36_clk_regs
+ sg13g2_dfrbpq_1
X_06914_ net3683 net2570 _02906_ _00697_ VPWR VGND sg13g2_a21o_1
X_07894_ i_exotiny._0021_\[2\] net876 _03228_ _03232_ VPWR VGND sg13g2_mux2_1
XFILLER_55_324 VPWR VGND sg13g2_decap_4
X_06845_ i_exotiny._0369_\[24\] net1188 _02858_ VPWR VGND sg13g2_nor2_1
X_06776_ _02800_ net1873 net1183 VPWR VGND sg13g2_nand2_1
X_08515_ net165 VGND VPWR net2275 i_exotiny._0043_\[3\] clknet_leaf_177_clk_regs sg13g2_dfrbpq_2
X_05727_ _02366_ net1105 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data[0]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_36_593 VPWR VGND sg13g2_fill_1
X_05658_ VGND VPWR net1063 _02314_ _00040_ _02312_ sg13g2_a21oi_1
X_08446_ net234 VGND VPWR _00520_ i_exotiny.i_wb_regs.spi_size_o\[0\] clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_2
X_08377_ net301 VGND VPWR net3267 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[15\]
+ clknet_leaf_134_clk_regs sg13g2_dfrbpq_1
X_04609_ _01371_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r VPWR VGND
+ sg13g2_inv_2
XFILLER_104_1000 VPWR VGND sg13g2_decap_8
X_05589_ net3390 _02263_ i_exotiny._1465_ VPWR VGND sg13g2_and2_1
X_07328_ _02992_ i_exotiny._0369_\[2\] i_exotiny._0369_\[3\] VPWR VGND sg13g2_nand2_2
XFILLER_87_1006 VPWR VGND sg13g2_decap_8
X_07259_ net2973 net2616 net1003 _00982_ VPWR VGND sg13g2_mux2_1
XFILLER_105_543 VPWR VGND sg13g2_decap_8
XFILLER_24_1001 VPWR VGND sg13g2_fill_1
X_08366__312 VPWR VGND net312 sg13g2_tiehi
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_104_93 VPWR VGND sg13g2_fill_1
XFILLER_15_777 VPWR VGND sg13g2_fill_1
XFILLER_6_420 VPWR VGND sg13g2_fill_1
XFILLER_7_954 VPWR VGND sg13g2_decap_8
XFILLER_50_7 VPWR VGND sg13g2_fill_2
X_08373__305 VPWR VGND net305 sg13g2_tiehi
X_09186__795 VPWR VGND net795 sg13g2_tiehi
Xclkbuf_5_28__f_clk_regs clknet_4_14_0_clk_regs clknet_5_28__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_09300__1117 VPWR VGND net1537 sg13g2_tiehi
XFILLER_29_4 VPWR VGND sg13g2_decap_4
X_04960_ _01690_ VPWR _01692_ VGND _01424_ _01691_ sg13g2_o21ai_1
XFILLER_93_942 VPWR VGND sg13g2_decap_8
X_08019__675 VPWR VGND net675 sg13g2_tiehi
XFILLER_92_452 VPWR VGND sg13g2_fill_1
X_04891_ _01623_ i_exotiny._0077_\[2\] VPWR VGND i_exotiny._0077_\[3\] sg13g2_nand2b_2
X_06630_ net1199 _02675_ _02676_ _00650_ VPWR VGND sg13g2_nor3_1
XFILLER_52_349 VPWR VGND sg13g2_fill_2
XFILLER_18_582 VPWR VGND sg13g2_fill_2
X_06561_ VGND VPWR _01394_ net1211 _00627_ _02630_ sg13g2_a21oi_1
X_09193__788 VPWR VGND net788 sg13g2_tiehi
X_08300_ net378 VGND VPWR _00381_ i_exotiny._0031_\[2\] clknet_leaf_72_clk_regs sg13g2_dfrbpq_2
X_06492_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[23\]
+ net2940 net1023 _00573_ VPWR VGND sg13g2_mux2_1
X_09280_ net61 VGND VPWR _01335_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[6\]
+ clknet_leaf_170_clk_regs sg13g2_dfrbpq_1
X_05512_ net1276 i_exotiny._0315_\[10\] _02204_ VPWR VGND sg13g2_nor2b_1
X_05443_ net1264 VPWR _02152_ VGND i_exotiny._1619_\[0\] _02138_ sg13g2_o21ai_1
X_08231_ net446 VGND VPWR net2665 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[30\]
+ clknet_leaf_151_clk_regs sg13g2_dfrbpq_1
X_08829__1159 VPWR VGND net1579 sg13g2_tiehi
X_05374_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set[0]
+ _02074_ _02095_ _02096_ VPWR VGND sg13g2_nor3_1
X_08162_ net516 VGND VPWR net2272 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[26\]
+ clknet_leaf_132_clk_regs sg13g2_dfrbpq_1
X_07113_ net1286 net1869 _00863_ VPWR VGND sg13g2_and2_1
X_08093_ net601 VGND VPWR net2478 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[30\]
+ clknet_leaf_85_clk_regs sg13g2_dfrbpq_1
X_08026__668 VPWR VGND net668 sg13g2_tiehi
XFILLER_106_307 VPWR VGND sg13g2_decap_8
X_07044_ net3194 net2920 net1017 _00805_ VPWR VGND sg13g2_mux2_1
XFILLER_88_703 VPWR VGND sg13g2_fill_2
XFILLER_87_224 VPWR VGND sg13g2_fill_1
XFILLER_87_213 VPWR VGND sg13g2_fill_1
X_08995_ net1407 VGND VPWR net3542 i_exotiny._1160_\[16\] clknet_leaf_18_clk_regs
+ sg13g2_dfrbpq_1
X_08072__622 VPWR VGND net622 sg13g2_tiehi
X_07946_ net90 VGND VPWR _00011_ i_exotiny._1711_ clknet_leaf_21_clk_regs sg13g2_dfrbpq_2
XFILLER_68_471 VPWR VGND sg13g2_decap_8
X_07877_ net2188 net2558 net980 _01344_ VPWR VGND sg13g2_mux2_1
XFILLER_18_57 VPWR VGND sg13g2_fill_1
XFILLER_70_102 VPWR VGND sg13g2_fill_1
X_06828_ net1170 VPWR _02844_ VGND net3600 net1185 sg13g2_o21ai_1
X_06759_ VGND VPWR _02786_ net1102 net1980 sg13g2_or2_1
XFILLER_34_89 VPWR VGND sg13g2_fill_2
X_08429_ net256 VGND VPWR net3325 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[28\]
+ clknet_leaf_91_clk_regs sg13g2_dfrbpq_1
Xclkload0 clkload0/Y clknet_5_2__leaf_clk_regs VPWR VGND sg13g2_inv_2
X_08402__283 VPWR VGND net283 sg13g2_tiehi
XFILLER_50_99 VPWR VGND sg13g2_fill_1
XFILLER_4_946 VPWR VGND sg13g2_decap_8
XFILLER_106_874 VPWR VGND sg13g2_decap_8
XFILLER_105_340 VPWR VGND sg13g2_decap_8
X_08872__1110 VPWR VGND net1530 sg13g2_tiehi
Xfanout1213 net1217 net1213 VPWR VGND sg13g2_buf_1
Xfanout1202 _01434_ net1202 VPWR VGND sg13g2_buf_1
Xfanout1246 net3807 net1246 VPWR VGND sg13g2_buf_1
Xfanout1235 net1237 net1235 VPWR VGND sg13g2_buf_8
Xfanout1224 _01382_ net1224 VPWR VGND sg13g2_buf_8
Xfanout1268 net3840 net1268 VPWR VGND sg13g2_buf_8
Xfanout1279 net1280 net1279 VPWR VGND sg13g2_buf_8
Xfanout1257 net3831 net1257 VPWR VGND sg13g2_buf_8
XFILLER_75_953 VPWR VGND sg13g2_fill_2
XFILLER_90_901 VPWR VGND sg13g2_fill_1
XFILLER_75_96 VPWR VGND sg13g2_fill_2
XFILLER_35_839 VPWR VGND sg13g2_fill_1
XFILLER_91_40 VPWR VGND sg13g2_fill_2
XFILLER_90_989 VPWR VGND sg13g2_decap_8
XFILLER_91_95 VPWR VGND sg13g2_fill_1
XFILLER_30_599 VPWR VGND sg13g2_fill_1
Xhold707 i_exotiny._0021_\[0\] VPWR VGND net2534 sg13g2_dlygate4sd3_1
Xhold718 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[9\]
+ VPWR VGND net2545 sg13g2_dlygate4sd3_1
Xhold729 _00818_ VPWR VGND net2556 sg13g2_dlygate4sd3_1
X_05090_ net1248 _01610_ _01821_ VPWR VGND sg13g2_nor2_1
Xhold1407 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[16\]
+ VPWR VGND net3234 sg13g2_dlygate4sd3_1
X_07800_ net2751 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[18\]
+ net893 _01279_ VPWR VGND sg13g2_mux2_1
X_08780_ net1628 VGND VPWR _00838_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[11\]
+ clknet_leaf_164_clk_regs sg13g2_dfrbpq_1
Xhold1429 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[6\]
+ VPWR VGND net3256 sg13g2_dlygate4sd3_1
Xhold1418 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[16\]
+ VPWR VGND net3245 sg13g2_dlygate4sd3_1
X_05992_ net3296 net3313 net1049 _00194_ VPWR VGND sg13g2_mux2_1
X_07731_ net3294 net886 _03199_ _03201_ VPWR VGND sg13g2_mux2_1
X_04943_ _01612_ _01673_ _01674_ _01675_ VPWR VGND sg13g2_nor3_1
X_07662_ net3145 _03192_ net897 _01166_ VPWR VGND sg13g2_mux2_1
X_04874_ _01605_ net1247 _01499_ _01606_ VPWR VGND sg13g2_a21o_1
X_07593_ net1179 VPWR _03167_ VGND net3642 _03165_ sg13g2_o21ai_1
XFILLER_53_647 VPWR VGND sg13g2_fill_1
XFILLER_52_124 VPWR VGND sg13g2_fill_1
X_06613_ net2864 net1160 _02665_ VPWR VGND sg13g2_nor2_1
XFILLER_37_187 VPWR VGND sg13g2_fill_1
XFILLER_52_146 VPWR VGND sg13g2_fill_2
X_06544_ net3239 _02624_ net929 _00616_ VPWR VGND sg13g2_mux2_1
XFILLER_40_308 VPWR VGND sg13g2_fill_1
X_06475_ net3482 i_exotiny._0041_\[2\] net1025 _00556_ VPWR VGND sg13g2_mux2_1
X_09263_ net235 VGND VPWR net2348 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[21\]
+ clknet_leaf_128_clk_regs sg13g2_dfrbpq_1
X_09194_ net787 VGND VPWR _01249_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[16\]
+ clknet_leaf_77_clk_regs sg13g2_dfrbpq_1
X_08950__1032 VPWR VGND net1452 sg13g2_tiehi
X_05426_ net1232 _02129_ _02134_ _02135_ VPWR VGND sg13g2_nor3_1
X_08214_ net463 VGND VPWR _00295_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[13\]
+ clknet_leaf_153_clk_regs sg13g2_dfrbpq_1
X_05357_ i_exotiny._2034_\[8\] _00022_ _02079_ VPWR VGND sg13g2_xor2_1
X_08145_ net540 VGND VPWR net2605 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[9\]
+ clknet_leaf_131_clk_regs sg13g2_dfrbpq_1
XFILLER_106_104 VPWR VGND sg13g2_decap_8
XFILLER_101_1025 VPWR VGND sg13g2_decap_4
X_08076_ net618 VGND VPWR net2171 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[13\]
+ clknet_leaf_92_clk_regs sg13g2_dfrbpq_1
X_08356__322 VPWR VGND net322 sg13g2_tiehi
X_05288_ _02012_ _01988_ _02013_ _02014_ VPWR VGND sg13g2_a21o_1
XFILLER_103_811 VPWR VGND sg13g2_decap_8
X_07027_ net3175 _02931_ net920 _00792_ VPWR VGND sg13g2_mux2_1
XFILLER_102_343 VPWR VGND sg13g2_decap_8
Xhold12 i_exotiny.i_wb_spi.state_r\[21\] VPWR VGND net1839 sg13g2_dlygate4sd3_1
Xhold23 _00871_ VPWR VGND net1850 sg13g2_dlygate4sd3_1
XFILLER_103_888 VPWR VGND sg13g2_decap_8
Xhold34 i_exotiny.i_wb_spi.state_r\[2\] VPWR VGND net1861 sg13g2_dlygate4sd3_1
Xhold56 i_exotiny.i_rstctl.cnt\[0\] VPWR VGND net1883 sg13g2_dlygate4sd3_1
Xhold45 i_exotiny._0369_\[26\] VPWR VGND net1872 sg13g2_dlygate4sd3_1
X_08978_ net1424 VGND VPWR _01036_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[3\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_2
XFILLER_75_249 VPWR VGND sg13g2_fill_2
Xhold78 i_exotiny.i_wb_spi.dat_rx_r\[12\] VPWR VGND net1905 sg13g2_dlygate4sd3_1
X_07929_ net719 VGND VPWR net1927 i_exotiny._1924_\[22\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
Xhold89 i_exotiny._1924_\[21\] VPWR VGND net1916 sg13g2_dlygate4sd3_1
Xhold1963 _01437_ VPWR VGND net3790 sg13g2_dlygate4sd3_1
Xhold1930 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[1\] VPWR VGND net3757
+ sg13g2_dlygate4sd3_1
Xhold67 _01495_ VPWR VGND net1894 sg13g2_dlygate4sd3_1
Xhold1941 i_exotiny._0369_\[4\] VPWR VGND net3768 sg13g2_dlygate4sd3_1
Xhold1952 _00512_ VPWR VGND net3779 sg13g2_dlygate4sd3_1
Xhold1974 i_exotiny._1615_\[3\] VPWR VGND net3801 sg13g2_dlygate4sd3_1
XFILLER_28_165 VPWR VGND sg13g2_fill_2
Xhold1996 _01072_ VPWR VGND net3823 sg13g2_dlygate4sd3_1
Xhold1985 i_exotiny._0077_\[1\] VPWR VGND net3812 sg13g2_dlygate4sd3_1
XFILLER_45_55 VPWR VGND sg13g2_fill_1
X_08363__315 VPWR VGND net315 sg13g2_tiehi
XFILLER_61_43 VPWR VGND sg13g2_fill_2
XFILLER_61_54 VPWR VGND sg13g2_fill_2
XFILLER_8_537 VPWR VGND sg13g2_fill_1
X_08770__1218 VPWR VGND net1638 sg13g2_tiehi
XFILLER_106_671 VPWR VGND sg13g2_decap_8
X_08370__308 VPWR VGND net308 sg13g2_tiehi
X_09183__798 VPWR VGND net798 sg13g2_tiehi
XFILLER_86_40 VPWR VGND sg13g2_fill_1
Xfanout1021 _02923_ net1021 VPWR VGND sg13g2_buf_8
Xfanout1010 _02948_ net1010 VPWR VGND sg13g2_buf_8
Xfanout1032 _02566_ net1032 VPWR VGND sg13g2_buf_8
Xfanout1065 net1066 net1065 VPWR VGND sg13g2_buf_8
Xfanout1054 net1055 net1054 VPWR VGND sg13g2_buf_8
Xfanout1043 net1045 net1043 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_129_clk_regs clknet_5_21__leaf_clk_regs clknet_leaf_129_clk_regs VPWR
+ VGND sg13g2_buf_8
Xfanout1098 net1099 net1098 VPWR VGND sg13g2_buf_1
Xfanout1087 net1091 net1087 VPWR VGND sg13g2_buf_1
Xfanout1076 _01526_ net1076 VPWR VGND sg13g2_buf_8
X_08016__678 VPWR VGND net678 sg13g2_tiehi
XFILLER_34_146 VPWR VGND sg13g2_fill_1
XFILLER_35_669 VPWR VGND sg13g2_fill_1
XFILLER_50_617 VPWR VGND sg13g2_decap_8
XFILLER_22_319 VPWR VGND sg13g2_fill_2
X_06260_ i_exotiny._0031_\[1\] net883 _02546_ _02549_ VPWR VGND sg13g2_mux2_1
X_08062__632 VPWR VGND net632 sg13g2_tiehi
X_09090__892 VPWR VGND net1312 sg13g2_tiehi
X_05211_ _01939_ _01772_ i_exotiny._0033_\[1\] _01758_ i_exotiny._0040_\[1\] VPWR
+ VGND sg13g2_a22oi_1
X_08746__1242 VPWR VGND net1662 sg13g2_tiehi
X_06191_ VGND VPWR net1140 _02540_ _02541_ net1166 sg13g2_a21oi_1
Xhold504 i_exotiny._1612_\[3\] VPWR VGND net2331 sg13g2_dlygate4sd3_1
Xhold515 _00584_ VPWR VGND net2342 sg13g2_dlygate4sd3_1
Xhold526 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[30\]
+ VPWR VGND net2353 sg13g2_dlygate4sd3_1
X_05142_ _01870_ _01845_ _01871_ _01872_ VPWR VGND sg13g2_a21o_1
Xhold537 _00581_ VPWR VGND net2364 sg13g2_dlygate4sd3_1
Xhold559 _00422_ VPWR VGND net2386 sg13g2_dlygate4sd3_1
Xhold548 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[20\]
+ VPWR VGND net2375 sg13g2_dlygate4sd3_1
X_05073_ _01764_ _01803_ _01755_ _01805_ VPWR VGND _01804_ sg13g2_nand4_1
XFILLER_103_129 VPWR VGND sg13g2_decap_8
X_08901_ net1501 VGND VPWR net3531 i_exotiny.i_wb_spi.dat_rx_r\[31\] clknet_leaf_19_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_98_853 VPWR VGND sg13g2_decap_8
XFILLER_97_352 VPWR VGND sg13g2_decap_8
X_08832_ net1576 VGND VPWR _00890_ i_exotiny.i_wb_spi.state_r\[31\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
Xhold1204 i_exotiny._0043_\[0\] VPWR VGND net3031 sg13g2_dlygate4sd3_1
Xhold1215 _00714_ VPWR VGND net3042 sg13g2_dlygate4sd3_1
XFILLER_100_847 VPWR VGND sg13g2_decap_8
Xhold1226 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[25\]
+ VPWR VGND net3053 sg13g2_dlygate4sd3_1
X_08763_ net1645 VGND VPWR net2314 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[26\]
+ clknet_leaf_84_clk_regs sg13g2_dfrbpq_1
XFILLER_73_709 VPWR VGND sg13g2_fill_1
Xhold1248 i_exotiny._0027_\[1\] VPWR VGND net3075 sg13g2_dlygate4sd3_1
Xhold1237 i_exotiny._0039_\[1\] VPWR VGND net3064 sg13g2_dlygate4sd3_1
XFILLER_39_953 VPWR VGND sg13g2_fill_2
X_05975_ net2946 net3532 net1049 _00177_ VPWR VGND sg13g2_mux2_1
X_07714_ net3198 net3176 net995 _01210_ VPWR VGND sg13g2_mux2_1
Xhold1259 _01163_ VPWR VGND net3086 sg13g2_dlygate4sd3_1
X_08968__1014 VPWR VGND net1434 sg13g2_tiehi
X_04926_ _01658_ _01652_ i_exotiny._0018_\[3\] _01649_ i_exotiny._0042_\[3\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_65_282 VPWR VGND sg13g2_fill_1
X_08694_ net1714 VGND VPWR _00752_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[21\]
+ clknet_leaf_116_clk_regs sg13g2_dfrbpq_1
XFILLER_25_124 VPWR VGND sg13g2_fill_2
XFILLER_80_252 VPWR VGND sg13g2_fill_2
X_04857_ _01592_ i_exotiny.i_wb_spi.cnt_presc_r\[5\] _01574_ VPWR VGND sg13g2_xnor2_1
X_07645_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[18\]
+ net2130 net897 _01153_ VPWR VGND sg13g2_mux2_1
X_07576_ _03155_ VPWR _03156_ VGND net3756 _03154_ sg13g2_o21ai_1
X_04788_ _01537_ net3713 _01538_ VPWR VGND sg13g2_xor2_1
XFILLER_90_1024 VPWR VGND sg13g2_decap_4
X_06527_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[16\]
+ net2701 net933 _00602_ VPWR VGND sg13g2_mux2_1
X_06458_ net3115 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[23\]
+ net935 _00545_ VPWR VGND sg13g2_mux2_1
X_09246_ net561 VGND VPWR _01301_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[4\]
+ clknet_leaf_126_clk_regs sg13g2_dfrbpq_1
X_05409_ i_exotiny._2034_\[7\] _02119_ _02121_ VPWR VGND sg13g2_and2_1
X_08499__181 VPWR VGND net181 sg13g2_tiehi
X_09177_ net805 VGND VPWR net1962 i_exotiny._1924_\[1\] clknet_leaf_30_clk_regs sg13g2_dfrbpq_1
X_06389_ _02576_ VPWR _00509_ VGND _01513_ _02131_ sg13g2_o21ai_1
X_08128_ net1178 VGND VPWR net1981 _00016_ clknet_leaf_36_clk_regs sg13g2_dfrbpq_1
X_08059_ net635 VGND VPWR net3121 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[28\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
Xoutput24 net24 uio_oe[6] VPWR VGND sg13g2_buf_1
Xoutput35 net35 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_89_875 VPWR VGND sg13g2_fill_2
XFILLER_1_768 VPWR VGND sg13g2_decap_8
XFILLER_48_205 VPWR VGND sg13g2_fill_1
XFILLER_88_396 VPWR VGND sg13g2_fill_1
Xhold1760 i_exotiny.i_wb_spi.dat_rx_r\[22\] VPWR VGND net3587 sg13g2_dlygate4sd3_1
XFILLER_63_219 VPWR VGND sg13g2_fill_1
Xhold1771 i_exotiny._1160_\[20\] VPWR VGND net3598 sg13g2_dlygate4sd3_1
Xhold1793 i_exotiny._1616_\[3\] VPWR VGND net3620 sg13g2_dlygate4sd3_1
Xhold1782 i_exotiny._1160_\[22\] VPWR VGND net3609 sg13g2_dlygate4sd3_1
X_08824__1164 VPWR VGND net1584 sg13g2_tiehi
XFILLER_32_628 VPWR VGND sg13g2_fill_1
XFILLER_44_488 VPWR VGND sg13g2_fill_1
XFILLER_31_127 VPWR VGND sg13g2_fill_1
XFILLER_8_323 VPWR VGND sg13g2_fill_1
X_09248__559 VPWR VGND net559 sg13g2_tiehi
XFILLER_98_127 VPWR VGND sg13g2_fill_2
XFILLER_67_525 VPWR VGND sg13g2_fill_2
XFILLER_95_856 VPWR VGND sg13g2_decap_8
XFILLER_94_344 VPWR VGND sg13g2_fill_2
XFILLER_94_333 VPWR VGND sg13g2_decap_8
XFILLER_94_355 VPWR VGND sg13g2_decap_4
X_05760_ _02391_ i_exotiny._2034_\[0\] net1127 VPWR VGND sg13g2_nand2_1
XFILLER_48_783 VPWR VGND sg13g2_fill_1
X_04711_ net1254 _01468_ _01469_ VPWR VGND sg13g2_nor2_1
X_07951__95 VPWR VGND net95 sg13g2_tiehi
X_05691_ net1123 net2046 _02339_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_97_clk_regs clknet_5_29__leaf_clk_regs clknet_leaf_97_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08346__332 VPWR VGND net332 sg13g2_tiehi
X_04642_ _01404_ i_exotiny._0369_\[6\] VPWR VGND sg13g2_inv_2
XFILLER_35_488 VPWR VGND sg13g2_fill_1
X_07430_ net1081 _03073_ _03074_ _03075_ VPWR VGND sg13g2_nor3_1
Xclkbuf_leaf_26_clk_regs clknet_5_9__leaf_clk_regs clknet_leaf_26_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07361_ net3647 net1213 _03021_ VPWR VGND sg13g2_and2_1
X_06312_ net3478 net3519 net1036 _00449_ VPWR VGND sg13g2_mux2_1
X_09100_ net1302 VGND VPWR net2237 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[20\]
+ clknet_leaf_142_clk_regs sg13g2_dfrbpq_1
X_07984__125 VPWR VGND net125 sg13g2_tiehi
X_07292_ net2127 net2295 net908 _01009_ VPWR VGND sg13g2_mux2_1
X_09031_ net1371 VGND VPWR _01089_ i_exotiny._0315_\[19\] clknet_leaf_180_clk_regs
+ sg13g2_dfrbpq_1
X_06243_ net2894 net3211 net1041 _00392_ VPWR VGND sg13g2_mux2_1
X_06174_ net3435 net3398 net953 _00336_ VPWR VGND sg13g2_mux2_1
Xhold301 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[5\]
+ VPWR VGND net2128 sg13g2_dlygate4sd3_1
Xhold312 _00475_ VPWR VGND net2139 sg13g2_dlygate4sd3_1
Xhold334 _00757_ VPWR VGND net2161 sg13g2_dlygate4sd3_1
Xhold323 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[29\]
+ VPWR VGND net2150 sg13g2_dlygate4sd3_1
X_05125_ _01852_ _01853_ _01850_ _01855_ VPWR VGND _01854_ sg13g2_nand4_1
Xhold378 _00892_ VPWR VGND net2205 sg13g2_dlygate4sd3_1
Xhold367 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[21\]
+ VPWR VGND net2194 sg13g2_dlygate4sd3_1
Xhold356 _01167_ VPWR VGND net2183 sg13g2_dlygate4sd3_1
Xhold345 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[30\]
+ VPWR VGND net2172 sg13g2_dlygate4sd3_1
X_08353__325 VPWR VGND net325 sg13g2_tiehi
Xhold389 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[31\]
+ VPWR VGND net2216 sg13g2_dlygate4sd3_1
X_05056_ net1236 _01757_ _01762_ _01788_ VPWR VGND sg13g2_nor3_2
XFILLER_98_672 VPWR VGND sg13g2_fill_2
X_08815_ net1593 VGND VPWR net1836 i_exotiny.i_wb_spi.state_r\[14\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
Xhold1001 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[9\]
+ VPWR VGND net2828 sg13g2_dlygate4sd3_1
Xhold1012 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[28\]
+ VPWR VGND net2839 sg13g2_dlygate4sd3_1
Xhold1023 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[21\]
+ VPWR VGND net2850 sg13g2_dlygate4sd3_1
Xhold1067 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[17\]
+ VPWR VGND net2894 sg13g2_dlygate4sd3_1
Xhold1056 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[17\]
+ VPWR VGND net2883 sg13g2_dlygate4sd3_1
Xhold1034 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[30\]
+ VPWR VGND net2861 sg13g2_dlygate4sd3_1
Xhold1045 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[12\]
+ VPWR VGND net2872 sg13g2_dlygate4sd3_1
X_08746_ net1662 VGND VPWR net1829 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[9\]
+ clknet_leaf_86_clk_regs sg13g2_dfrbpq_1
X_05958_ net2456 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[27\]
+ net969 _00167_ VPWR VGND sg13g2_mux2_1
Xhold1089 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[16\]
+ VPWR VGND net2916 sg13g2_dlygate4sd3_1
Xhold1078 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[4\]
+ VPWR VGND net2905 sg13g2_dlygate4sd3_1
XFILLER_53_230 VPWR VGND sg13g2_fill_1
X_08677_ net1731 VGND VPWR net3310 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[4\]
+ clknet_leaf_102_clk_regs sg13g2_dfrbpq_1
X_05889_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[0\] _02417_ _02474_
+ VPWR VGND sg13g2_nor2b_1
X_04909_ net1222 _01613_ _01640_ _01641_ VPWR VGND sg13g2_nor3_2
XFILLER_54_775 VPWR VGND sg13g2_fill_1
X_07628_ i_exotiny._0024_\[1\] net2186 net898 _01136_ VPWR VGND sg13g2_mux2_1
XFILLER_53_285 VPWR VGND sg13g2_fill_1
X_07559_ VGND VPWR net1970 _03142_ _01111_ _03144_ sg13g2_a21oi_1
X_08360__318 VPWR VGND net318 sg13g2_tiehi
X_09229_ net750 VGND VPWR net2346 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[19\]
+ clknet_leaf_134_clk_regs sg13g2_dfrbpq_1
XFILLER_42_89 VPWR VGND sg13g2_fill_1
XFILLER_10_889 VPWR VGND sg13g2_fill_1
Xhold890 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[27\]
+ VPWR VGND net2717 sg13g2_dlygate4sd3_1
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_104_972 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_fill_1
XFILLER_103_493 VPWR VGND sg13g2_decap_8
X_08052__642 VPWR VGND net642 sg13g2_tiehi
Xhold1590 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[4\]
+ VPWR VGND net3417 sg13g2_dlygate4sd3_1
XFILLER_40_491 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_144_clk_regs clknet_5_17__leaf_clk_regs clknet_leaf_144_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_5_882 VPWR VGND sg13g2_decap_8
XFILLER_102_909 VPWR VGND sg13g2_decap_8
XFILLER_99_458 VPWR VGND sg13g2_decap_8
XFILLER_87_609 VPWR VGND sg13g2_fill_1
XFILLER_101_408 VPWR VGND sg13g2_decap_8
X_06930_ net2783 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[14\]
+ net925 _00709_ VPWR VGND sg13g2_mux2_1
X_08600_ net1796 VGND VPWR _00672_ i_exotiny._1615_\[0\] clknet_leaf_58_clk_regs sg13g2_dfrbpq_2
X_08696__1292 VPWR VGND net1712 sg13g2_tiehi
X_06861_ net3614 net1095 _02872_ VPWR VGND sg13g2_nor2_1
X_08489__191 VPWR VGND net191 sg13g2_tiehi
X_05812_ net2085 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[4\]
+ net1055 _00084_ VPWR VGND sg13g2_mux2_1
X_06792_ VGND VPWR net3711 net1133 _02814_ _02813_ sg13g2_a21oi_1
X_05743_ _02373_ _02376_ _02379_ VPWR VGND sg13g2_nor2_1
X_08531_ net149 VGND VPWR _00605_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[19\]
+ clknet_leaf_182_clk_regs sg13g2_dfrbpq_1
X_05674_ VGND VPWR net1062 _02326_ _00044_ _02324_ sg13g2_a21oi_1
X_08462_ net218 VGND VPWR net2649 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[14\]
+ clknet_leaf_114_clk_regs sg13g2_dfrbpq_1
XFILLER_51_734 VPWR VGND sg13g2_fill_1
XFILLER_50_222 VPWR VGND sg13g2_fill_1
X_08591__1385 VPWR VGND net1805 sg13g2_tiehi
XFILLER_23_447 VPWR VGND sg13g2_fill_2
X_07413_ VGND VPWR i_exotiny._0369_\[15\] net1147 _03062_ _03052_ sg13g2_a21oi_1
X_04625_ VPWR _01387_ net3789 VGND sg13g2_inv_1
X_08393_ net533 VGND VPWR _00474_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[31\]
+ clknet_leaf_141_clk_regs sg13g2_dfrbpq_1
X_07344_ VGND VPWR net1078 _03006_ _01033_ _03007_ sg13g2_a21oi_1
X_07275_ i_exotiny._0042_\[0\] net2438 net910 _00992_ VPWR VGND sg13g2_mux2_1
X_06226_ i_exotiny._0033_\[3\] net874 _02540_ _02545_ VPWR VGND sg13g2_mux2_1
X_09014_ net1388 VGND VPWR net3823 i_exotiny._0315_\[2\] clknet_leaf_11_clk_regs sg13g2_dfrbpq_2
X_08496__184 VPWR VGND net184 sg13g2_tiehi
X_06157_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[5\]
+ net3277 net951 _00319_ VPWR VGND sg13g2_mux2_1
Xhold153 i_exotiny._1612_\[2\] VPWR VGND net1980 sg13g2_dlygate4sd3_1
Xhold142 _00936_ VPWR VGND net1969 sg13g2_dlygate4sd3_1
Xhold120 i_exotiny._1924_\[19\] VPWR VGND net1947 sg13g2_dlygate4sd3_1
Xhold131 _00045_ VPWR VGND net1958 sg13g2_dlygate4sd3_1
XFILLER_105_769 VPWR VGND sg13g2_decap_8
Xhold164 i_exotiny.i_wb_spi.cnt_hbit_r\[3\] VPWR VGND net1991 sg13g2_dlygate4sd3_1
X_06088_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[14\]
+ net2619 net958 _00264_ VPWR VGND sg13g2_mux2_1
Xhold186 _00216_ VPWR VGND net2013 sg13g2_dlygate4sd3_1
Xhold175 i_exotiny._0314_\[29\] VPWR VGND net2002 sg13g2_dlygate4sd3_1
X_05108_ VGND VPWR _01838_ _01742_ _01720_ sg13g2_or2_1
XFILLER_104_257 VPWR VGND sg13g2_decap_8
Xhold197 i_exotiny._0315_\[31\] VPWR VGND net2024 sg13g2_dlygate4sd3_1
X_05039_ net1235 _01754_ _01762_ _01771_ VPWR VGND sg13g2_nor3_2
XFILLER_101_920 VPWR VGND sg13g2_decap_8
XFILLER_86_620 VPWR VGND sg13g2_fill_1
XFILLER_100_430 VPWR VGND sg13g2_decap_8
XFILLER_58_355 VPWR VGND sg13g2_fill_1
XFILLER_101_997 VPWR VGND sg13g2_decap_8
XFILLER_27_731 VPWR VGND sg13g2_fill_2
X_08729_ net1679 VGND VPWR net2084 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[24\]
+ clknet_leaf_119_clk_regs sg13g2_dfrbpq_1
XFILLER_39_591 VPWR VGND sg13g2_fill_1
XFILLER_27_775 VPWR VGND sg13g2_fill_2
XFILLER_27_797 VPWR VGND sg13g2_fill_1
XFILLER_41_200 VPWR VGND sg13g2_fill_1
XFILLER_6_602 VPWR VGND sg13g2_fill_1
Xclkbuf_5_27__f_clk_regs clknet_4_13_0_clk_regs clknet_5_27__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_2_852 VPWR VGND sg13g2_decap_8
X_08336__342 VPWR VGND net342 sg13g2_tiehi
XFILLER_77_642 VPWR VGND sg13g2_fill_1
XFILLER_103_290 VPWR VGND sg13g2_decap_8
XFILLER_49_344 VPWR VGND sg13g2_fill_2
XFILLER_45_572 VPWR VGND sg13g2_decap_8
XFILLER_33_723 VPWR VGND sg13g2_fill_1
XFILLER_45_583 VPWR VGND sg13g2_fill_2
X_08343__335 VPWR VGND net335 sg13g2_tiehi
XFILLER_60_542 VPWR VGND sg13g2_fill_1
X_05390_ i_exotiny._2034_\[0\] net1112 i_exotiny._2043_\[0\] VPWR VGND sg13g2_nor2_1
XFILLER_14_981 VPWR VGND sg13g2_decap_8
XFILLER_20_439 VPWR VGND sg13g2_fill_1
X_07060_ net2313 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[26\]
+ net1017 _00821_ VPWR VGND sg13g2_mux2_1
X_06011_ VGND VPWR net3142 net1105 _00208_ _02499_ sg13g2_a21oi_1
X_09048__804 VPWR VGND net804 sg13g2_tiehi
XFILLER_101_205 VPWR VGND sg13g2_decap_8
XFILLER_99_255 VPWR VGND sg13g2_decap_8
X_07962_ net1176 VGND VPWR net3529 i_exotiny.i_wdg_top.o_wb_dat\[3\] clknet_leaf_37_clk_regs
+ sg13g2_dfrbpq_2
X_08350__328 VPWR VGND net328 sg13g2_tiehi
X_08783__1205 VPWR VGND net1625 sg13g2_tiehi
XFILLER_96_984 VPWR VGND sg13g2_decap_8
X_06913_ _01389_ net3682 net1883 _02913_ VPWR VGND _02912_ sg13g2_nand4_1
X_07893_ net3097 _03231_ net978 _01358_ VPWR VGND sg13g2_mux2_1
XFILLER_95_472 VPWR VGND sg13g2_fill_2
X_06844_ VGND VPWR net1097 _02856_ _00683_ _02857_ sg13g2_a21oi_1
Xclkbuf_leaf_41_clk_regs clknet_5_10__leaf_clk_regs clknet_leaf_41_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06775_ VGND VPWR net1100 _02798_ _00672_ _02799_ sg13g2_a21oi_1
X_08514_ net166 VGND VPWR net3095 i_exotiny._0043_\[2\] clknet_leaf_183_clk_regs sg13g2_dfrbpq_2
X_05726_ VGND VPWR net1058 _02364_ _00057_ _02365_ sg13g2_a21oi_1
X_05657_ VGND VPWR i_exotiny._1614_\[2\] net1122 _02314_ _02313_ sg13g2_a21oi_1
X_08445_ net236 VGND VPWR _00519_ i_exotiny.i_wb_qspi_mem.crm_r clknet_leaf_16_clk_regs
+ sg13g2_dfrbpq_2
X_08376_ net302 VGND VPWR net3258 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[14\]
+ clknet_leaf_137_clk_regs sg13g2_dfrbpq_1
X_04608_ _01370_ net2886 VPWR VGND sg13g2_inv_2
X_05588_ _02262_ i_exotiny._0314_\[2\] _02263_ VPWR VGND sg13g2_nor2b_1
X_07327_ _02991_ net1208 _02989_ VPWR VGND sg13g2_nand2_2
X_07258_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[25\]
+ net2713 net1005 _00981_ VPWR VGND sg13g2_mux2_1
X_08042__652 VPWR VGND net652 sg13g2_tiehi
X_06209_ net2369 net2643 net946 _00364_ VPWR VGND sg13g2_mux2_1
X_07189_ net1281 VPWR _02959_ VGND net3744 _02956_ sg13g2_o21ai_1
XFILLER_105_522 VPWR VGND sg13g2_decap_8
XFILLER_105_599 VPWR VGND sg13g2_decap_8
XFILLER_48_33 VPWR VGND sg13g2_fill_1
XFILLER_101_750 VPWR VGND sg13g2_decap_8
XFILLER_47_804 VPWR VGND sg13g2_fill_2
XFILLER_101_794 VPWR VGND sg13g2_decap_8
XFILLER_64_87 VPWR VGND sg13g2_fill_1
XFILLER_61_328 VPWR VGND sg13g2_fill_2
XFILLER_54_380 VPWR VGND sg13g2_fill_2
XFILLER_11_995 VPWR VGND sg13g2_decap_8
XFILLER_7_933 VPWR VGND sg13g2_decap_8
XFILLER_31_1028 VPWR VGND sg13g2_fill_1
X_08904__1078 VPWR VGND net1498 sg13g2_tiehi
X_08579__1404 VPWR VGND net1824 sg13g2_tiehi
XFILLER_93_921 VPWR VGND sg13g2_decap_8
X_04890_ i_exotiny._0077_\[2\] i_exotiny._0077_\[3\] net1256 _01622_ VGND VPWR _01620_
+ sg13g2_nor4_2
XFILLER_93_998 VPWR VGND sg13g2_decap_8
X_08486__194 VPWR VGND net194 sg13g2_tiehi
XFILLER_46_870 VPWR VGND sg13g2_fill_2
X_06560_ net3505 _01504_ _02630_ VPWR VGND sg13g2_nor2_1
X_06491_ net3012 net3021 net1027 _00572_ VPWR VGND sg13g2_mux2_1
X_05511_ _02203_ net3307 net1069 VPWR VGND sg13g2_nand2_1
X_05442_ _02141_ _02147_ _02139_ _02151_ VPWR VGND _02150_ sg13g2_nand4_1
X_08230_ net447 VGND VPWR net2683 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[29\]
+ clknet_leaf_153_clk_regs sg13g2_dfrbpq_1
X_05373_ net1832 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.genblk7.g_value.r_value[0]
+ _02095_ VPWR VGND sg13g2_nor2b_1
X_08161_ net517 VGND VPWR _00242_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[25\]
+ clknet_leaf_133_clk_regs sg13g2_dfrbpq_1
X_07112_ net1288 net1851 _00862_ VPWR VGND sg13g2_and2_1
X_08092_ net602 VGND VPWR net2773 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[29\]
+ clknet_leaf_86_clk_regs sg13g2_dfrbpq_1
X_07043_ net1828 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[9\]
+ net1015 _00804_ VPWR VGND sg13g2_mux2_1
Xclkload40 clknet_leaf_82_clk_regs clkload40/X VPWR VGND sg13g2_buf_8
X_08493__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_102_525 VPWR VGND sg13g2_decap_4
X_08994_ net1408 VGND VPWR net2021 i_exotiny._1160_\[15\] clknet_leaf_162_clk_regs
+ sg13g2_dfrbpq_1
X_07945_ net89 VGND VPWR net3653 i_exotiny._1757_ clknet_leaf_10_clk_regs sg13g2_dfrbpq_2
XFILLER_96_792 VPWR VGND sg13g2_fill_2
X_07876_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[14\]
+ net3250 net981 _01343_ VPWR VGND sg13g2_mux2_1
XFILLER_29_848 VPWR VGND sg13g2_fill_2
X_06827_ net2125 net1188 _02843_ VPWR VGND sg13g2_nor2_1
X_06758_ VPWR VGND net3656 _02784_ net3821 net3835 _02785_ net1182 sg13g2_a221oi_1
X_05709_ VGND VPWR i_exotiny._1619_\[3\] net1115 _02353_ _02352_ sg13g2_a21oi_1
X_09239__697 VPWR VGND net697 sg13g2_tiehi
X_08326__352 VPWR VGND net352 sg13g2_tiehi
X_08428_ net257 VGND VPWR _00502_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[27\]
+ clknet_leaf_96_clk_regs sg13g2_dfrbpq_1
X_06689_ _02726_ _02725_ i_exotiny.gpo\[0\] _02722_ net1116 VPWR VGND sg13g2_a22oi_1
XFILLER_54_1028 VPWR VGND sg13g2_fill_1
XFILLER_51_361 VPWR VGND sg13g2_fill_1
X_07900__46 VPWR VGND net46 sg13g2_tiehi
X_08359_ net319 VGND VPWR net2425 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[29\]
+ clknet_leaf_94_clk_regs sg13g2_dfrbpq_1
XFILLER_50_23 VPWR VGND sg13g2_fill_2
Xclkload1 clknet_5_7__leaf_clk_regs clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_4_925 VPWR VGND sg13g2_decap_8
XFILLER_106_853 VPWR VGND sg13g2_decap_8
XFILLER_79_704 VPWR VGND sg13g2_fill_1
XFILLER_105_396 VPWR VGND sg13g2_decap_8
Xfanout1203 i_exotiny.i_wdg_top.cntr_inst.rst_n_sync net1203 VPWR VGND sg13g2_buf_8
Xfanout1214 net1217 net1214 VPWR VGND sg13g2_buf_8
X_08333__345 VPWR VGND net345 sg13g2_tiehi
Xfanout1225 net1226 net1225 VPWR VGND sg13g2_buf_8
Xfanout1247 i_exotiny._0590_ net1247 VPWR VGND sg13g2_buf_8
Xfanout1236 net1237 net1236 VPWR VGND sg13g2_buf_8
XFILLER_75_932 VPWR VGND sg13g2_fill_2
Xfanout1269 net3840 net1269 VPWR VGND sg13g2_buf_1
Xfanout1258 net1259 net1258 VPWR VGND sg13g2_buf_8
XFILLER_75_42 VPWR VGND sg13g2_fill_2
XFILLER_19_325 VPWR VGND sg13g2_fill_2
XFILLER_19_347 VPWR VGND sg13g2_fill_1
XFILLER_90_968 VPWR VGND sg13g2_decap_8
XFILLER_30_523 VPWR VGND sg13g2_fill_2
X_08340__338 VPWR VGND net338 sg13g2_tiehi
Xhold719 _01208_ VPWR VGND net2546 sg13g2_dlygate4sd3_1
Xhold708 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[5\]
+ VPWR VGND net2535 sg13g2_dlygate4sd3_1
XFILLER_3_991 VPWR VGND sg13g2_decap_8
XFILLER_69_258 VPWR VGND sg13g2_fill_1
Xhold1408 i_exotiny.i_wdg_top.clk_div_inst.cnt\[13\] VPWR VGND net3235 sg13g2_dlygate4sd3_1
Xhold1419 _00326_ VPWR VGND net3246 sg13g2_dlygate4sd3_1
XFILLER_66_910 VPWR VGND sg13g2_fill_2
X_05991_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[17\]
+ net3487 net1050 _00193_ VPWR VGND sg13g2_mux2_1
X_07730_ net2547 net2387 net993 _01226_ VPWR VGND sg13g2_mux2_1
XFILLER_66_965 VPWR VGND sg13g2_fill_1
X_04942_ i_exotiny._0036_\[3\] _01644_ _01674_ VPWR VGND sg13g2_nor2_1
X_07661_ i_exotiny._0024_\[3\] net873 _03187_ _03192_ VPWR VGND sg13g2_mux2_1
X_04873_ net1242 _01604_ _01605_ VPWR VGND sg13g2_nor2_1
X_07592_ net3642 _03165_ _03166_ VPWR VGND sg13g2_and2_1
X_08032__662 VPWR VGND net662 sg13g2_tiehi
XFILLER_77_1028 VPWR VGND sg13g2_fill_1
X_06612_ net1194 _02663_ _02664_ _00644_ VPWR VGND sg13g2_nor3_1
XFILLER_25_339 VPWR VGND sg13g2_fill_1
X_06543_ i_exotiny._0043_\[2\] net876 _02620_ _02624_ VPWR VGND sg13g2_mux2_1
XFILLER_21_501 VPWR VGND sg13g2_fill_1
XFILLER_33_361 VPWR VGND sg13g2_fill_2
XFILLER_34_873 VPWR VGND sg13g2_fill_1
X_06474_ net2983 net3133 net1024 _00555_ VPWR VGND sg13g2_mux2_1
X_09262_ net237 VGND VPWR net2470 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[20\]
+ clknet_leaf_127_clk_regs sg13g2_dfrbpq_1
X_09193_ net788 VGND VPWR _01248_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[15\]
+ clknet_leaf_77_clk_regs sg13g2_dfrbpq_1
X_05425_ _02134_ _01383_ _02131_ VPWR VGND sg13g2_xnor2_1
X_08213_ net464 VGND VPWR net3015 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[12\]
+ clknet_leaf_149_clk_regs sg13g2_dfrbpq_1
XFILLER_14_1001 VPWR VGND sg13g2_fill_2
XFILLER_14_1012 VPWR VGND sg13g2_decap_8
XFILLER_21_567 VPWR VGND sg13g2_fill_1
XFILLER_101_1004 VPWR VGND sg13g2_decap_8
X_05356_ _02078_ _00018_ i_exotiny._2034_\[4\] VPWR VGND sg13g2_xnor2_1
X_08144_ net541 VGND VPWR _00225_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[8\]
+ clknet_leaf_131_clk_regs sg13g2_dfrbpq_1
XFILLER_105_9 VPWR VGND sg13g2_fill_1
X_08075_ net619 VGND VPWR net2793 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[12\]
+ clknet_leaf_89_clk_regs sg13g2_dfrbpq_1
X_05287_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[0\] net1107
+ _02013_ VPWR VGND sg13g2_and2_1
X_07026_ net3202 net884 _02928_ _02931_ VPWR VGND sg13g2_mux2_1
XFILLER_103_867 VPWR VGND sg13g2_decap_8
XFILLER_102_322 VPWR VGND sg13g2_decap_8
Xhold13 i_exotiny.i_wb_spi.cnt_presc_r\[0\] VPWR VGND net1840 sg13g2_dlygate4sd3_1
Xhold35 i_exotiny.i_wb_spi.state_r\[24\] VPWR VGND net1862 sg13g2_dlygate4sd3_1
Xhold24 i_exotiny.i_wb_spi.state_r\[3\] VPWR VGND net1851 sg13g2_dlygate4sd3_1
Xhold46 i_exotiny.i_wdg_top.o_wb_dat\[13\] VPWR VGND net1873 sg13g2_dlygate4sd3_1
Xhold1920 i_exotiny._1619_\[3\] VPWR VGND net3747 sg13g2_dlygate4sd3_1
X_08977_ net1425 VGND VPWR _01035_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[2\]
+ clknet_leaf_165_clk_regs sg13g2_dfrbpq_2
XFILLER_102_399 VPWR VGND sg13g2_decap_8
Xhold1953 i_exotiny.i_wdg_top.do_cnt VPWR VGND net3780 sg13g2_dlygate4sd3_1
Xhold57 _01105_ VPWR VGND net1884 sg13g2_dlygate4sd3_1
Xhold79 _00941_ VPWR VGND net1906 sg13g2_dlygate4sd3_1
Xhold68 i_exotiny._1924_\[7\] VPWR VGND net1895 sg13g2_dlygate4sd3_1
X_07928_ net720 VGND VPWR net1917 i_exotiny._1924_\[21\] clknet_leaf_26_clk_regs sg13g2_dfrbpq_1
XFILLER_56_431 VPWR VGND sg13g2_fill_2
Xhold1931 _00619_ VPWR VGND net3758 sg13g2_dlygate4sd3_1
X_08860__1126 VPWR VGND net1546 sg13g2_tiehi
Xhold1942 _01026_ VPWR VGND net3769 sg13g2_dlygate4sd3_1
Xhold1964 i_exotiny.i_wdg_top.o_wb_dat\[9\] VPWR VGND net3791 sg13g2_dlygate4sd3_1
XFILLER_28_144 VPWR VGND sg13g2_fill_1
X_07859_ _03227_ net2267 net983 _01328_ VPWR VGND sg13g2_mux2_1
Xhold1986 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[5\] VPWR
+ VGND net3813 sg13g2_dlygate4sd3_1
Xhold1975 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[3\]
+ VPWR VGND net3802 sg13g2_dlygate4sd3_1
Xhold1997 i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[0\] VPWR VGND net3824 sg13g2_dlygate4sd3_1
XFILLER_25_862 VPWR VGND sg13g2_fill_2
X_08009__686 VPWR VGND net686 sg13g2_tiehi
XFILLER_4_700 VPWR VGND sg13g2_fill_1
Xclkbuf_4_8_0_clk_regs clknet_0_clk_regs clknet_4_8_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_106_650 VPWR VGND sg13g2_decap_8
XFILLER_3_243 VPWR VGND sg13g2_fill_2
XFILLER_4_799 VPWR VGND sg13g2_decap_8
XFILLER_105_193 VPWR VGND sg13g2_decap_8
XFILLER_79_545 VPWR VGND sg13g2_decap_8
Xfanout1022 _02923_ net1022 VPWR VGND sg13g2_buf_2
XFILLER_10_92 VPWR VGND sg13g2_fill_1
Xfanout1011 net1012 net1011 VPWR VGND sg13g2_buf_8
Xfanout1000 net1002 net1000 VPWR VGND sg13g2_buf_8
Xfanout1055 _02424_ net1055 VPWR VGND sg13g2_buf_8
Xfanout1033 net1034 net1033 VPWR VGND sg13g2_buf_8
Xfanout1044 net1045 net1044 VPWR VGND sg13g2_buf_1
X_09079__903 VPWR VGND net1323 sg13g2_tiehi
Xfanout1066 net1067 net1066 VPWR VGND sg13g2_buf_8
Xfanout1088 net1090 net1088 VPWR VGND sg13g2_buf_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
Xfanout1077 _02991_ net1077 VPWR VGND sg13g2_buf_8
Xfanout1099 net1100 net1099 VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_169_clk_regs clknet_5_5__leaf_clk_regs clknet_leaf_169_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_19_166 VPWR VGND sg13g2_fill_1
X_09257__550 VPWR VGND net550 sg13g2_tiehi
XFILLER_47_497 VPWR VGND sg13g2_fill_2
X_08483__197 VPWR VGND net197 sg13g2_tiehi
XFILLER_96_5 VPWR VGND sg13g2_fill_2
X_06190_ _02509_ _02532_ _02540_ VPWR VGND sg13g2_nor2_2
X_05210_ VPWR VGND i_exotiny._0042_\[1\] _01937_ _01784_ i_exotiny._0027_\[1\] _01938_
+ _01765_ sg13g2_a221oi_1
X_05141_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[2\] net1108
+ _01871_ VPWR VGND sg13g2_and2_1
Xhold505 _00210_ VPWR VGND net2332 sg13g2_dlygate4sd3_1
Xhold516 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[20\]
+ VPWR VGND net2343 sg13g2_dlygate4sd3_1
Xhold527 _00473_ VPWR VGND net2354 sg13g2_dlygate4sd3_1
Xhold549 _00367_ VPWR VGND net2376 sg13g2_dlygate4sd3_1
Xhold538 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[9\]
+ VPWR VGND net2365 sg13g2_dlygate4sd3_1
X_05072_ _01804_ _01792_ i_exotiny._0038_\[3\] _01771_ i_exotiny._0016_\[3\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_103_108 VPWR VGND sg13g2_fill_1
XFILLER_98_832 VPWR VGND sg13g2_decap_8
XFILLER_83_1021 VPWR VGND sg13g2_decap_8
X_08900_ net1502 VGND VPWR net3583 i_exotiny.i_wb_spi.dat_rx_r\[30\] clknet_leaf_21_clk_regs
+ sg13g2_dfrbpq_1
X_08831_ net1577 VGND VPWR _00889_ i_exotiny.i_wb_spi.state_r\[30\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_97_331 VPWR VGND sg13g2_decap_8
X_08641__1336 VPWR VGND net1756 sg13g2_tiehi
XFILLER_44_1027 VPWR VGND sg13g2_fill_2
XFILLER_100_826 VPWR VGND sg13g2_decap_8
X_08316__362 VPWR VGND net362 sg13g2_tiehi
Xhold1205 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[20\]
+ VPWR VGND net3032 sg13g2_dlygate4sd3_1
Xhold1216 i_exotiny._0029_\[2\] VPWR VGND net3043 sg13g2_dlygate4sd3_1
Xhold1238 i_exotiny._0017_\[3\] VPWR VGND net3065 sg13g2_dlygate4sd3_1
X_08762_ net1646 VGND VPWR net2807 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[25\]
+ clknet_leaf_87_clk_regs sg13g2_dfrbpq_1
XFILLER_57_228 VPWR VGND sg13g2_fill_2
Xhold1227 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[17\]
+ VPWR VGND net3054 sg13g2_dlygate4sd3_1
Xhold1249 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[12\]
+ VPWR VGND net3076 sg13g2_dlygate4sd3_1
X_05974_ i_exotiny._0013_\[0\] net3417 net1051 _00176_ VPWR VGND sg13g2_mux2_1
X_08693_ net1715 VGND VPWR net2909 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[20\]
+ clknet_leaf_102_clk_regs sg13g2_dfrbpq_1
X_07713_ net3271 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[10\]
+ net995 _01209_ VPWR VGND sg13g2_mux2_1
X_04925_ _01657_ _01650_ i_exotiny._0016_\[3\] _01625_ i_exotiny._0030_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_07644_ net3311 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[21\]
+ net898 _01152_ VPWR VGND sg13g2_mux2_1
XFILLER_25_114 VPWR VGND sg13g2_fill_1
X_04856_ VGND VPWR net1072 _01590_ i_exotiny._1902_\[4\] _01591_ sg13g2_a21oi_1
XFILLER_54_979 VPWR VGND sg13g2_fill_1
XFILLER_53_467 VPWR VGND sg13g2_fill_1
X_07575_ VGND VPWR net3756 _03154_ _03155_ net1204 sg13g2_a21oi_1
XFILLER_90_1003 VPWR VGND sg13g2_decap_8
X_04787_ VGND VPWR net1243 _01437_ _01537_ net1273 sg13g2_a21oi_1
X_06526_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[15\]
+ net2224 net930 _00601_ VPWR VGND sg13g2_mux2_1
X_06457_ net3342 net2667 net937 _00544_ VPWR VGND sg13g2_mux2_1
XFILLER_21_364 VPWR VGND sg13g2_fill_2
X_09245_ net562 VGND VPWR net2308 i_exotiny._0022_\[3\] clknet_leaf_131_clk_regs sg13g2_dfrbpq_2
X_05408_ i_exotiny._2034_\[7\] _02119_ _02120_ VPWR VGND sg13g2_nor2_1
X_08323__355 VPWR VGND net355 sg13g2_tiehi
X_09176_ net806 VGND VPWR net3806 i_exotiny.i_wb_spi.sck_r clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_1
X_06388_ VGND VPWR net3764 _02180_ _02576_ net1225 sg13g2_a21oi_1
XFILLER_31_47 VPWR VGND sg13g2_decap_8
X_08127_ net1176 VGND VPWR net3143 _00015_ clknet_leaf_37_clk_regs sg13g2_dfrbpq_1
X_05339_ _01828_ _02062_ _02063_ VPWR VGND sg13g2_nor2b_1
X_08058_ net636 VGND VPWR _00139_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[27\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
Xoutput25 net25 uio_oe[7] VPWR VGND sg13g2_buf_1
Xoutput36 net36 uo_out[2] VPWR VGND sg13g2_buf_1
X_07009_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[13\]
+ net2075 net921 _00776_ VPWR VGND sg13g2_mux2_1
XFILLER_88_320 VPWR VGND sg13g2_fill_2
XFILLER_1_747 VPWR VGND sg13g2_decap_8
XFILLER_102_196 VPWR VGND sg13g2_decap_8
X_08330__348 VPWR VGND net348 sg13g2_tiehi
Xhold1761 _00951_ VPWR VGND net3588 sg13g2_dlygate4sd3_1
Xhold1750 _00930_ VPWR VGND net3577 sg13g2_dlygate4sd3_1
Xhold1794 _00687_ VPWR VGND net3621 sg13g2_dlygate4sd3_1
Xhold1783 i_exotiny._0314_\[22\] VPWR VGND net3610 sg13g2_dlygate4sd3_1
Xhold1772 _01057_ VPWR VGND net3599 sg13g2_dlygate4sd3_1
XFILLER_16_125 VPWR VGND sg13g2_fill_2
XFILLER_44_434 VPWR VGND sg13g2_fill_1
XFILLER_13_821 VPWR VGND sg13g2_fill_1
XFILLER_4_530 VPWR VGND sg13g2_fill_2
X_08022__672 VPWR VGND net672 sg13g2_tiehi
XFILLER_94_312 VPWR VGND sg13g2_decap_8
XFILLER_0_791 VPWR VGND sg13g2_decap_8
XFILLER_48_773 VPWR VGND sg13g2_fill_1
X_04710_ _01468_ net1243 _01421_ VPWR VGND sg13g2_nand2_1
X_05690_ VGND VPWR net1062 _02338_ _00048_ _02336_ sg13g2_a21oi_1
XFILLER_62_242 VPWR VGND sg13g2_fill_1
XFILLER_63_776 VPWR VGND sg13g2_fill_1
X_04641_ _01403_ net3768 VPWR VGND sg13g2_inv_2
X_07360_ net3803 VPWR _01036_ VGND net1079 _03019_ sg13g2_o21ai_1
XFILLER_50_459 VPWR VGND sg13g2_fill_1
X_06311_ net2538 net2465 net1033 _00448_ VPWR VGND sg13g2_mux2_1
X_07291_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[16\]
+ net2245 net910 _01008_ VPWR VGND sg13g2_mux2_1
X_08659__1318 VPWR VGND net1738 sg13g2_tiehi
X_09030_ net1372 VGND VPWR net3550 i_exotiny._0315_\[18\] clknet_leaf_167_clk_regs
+ sg13g2_dfrbpq_1
X_06242_ net2621 net3213 net1041 _00391_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_66_clk_regs clknet_5_24__leaf_clk_regs clknet_leaf_66_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06173_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[21\]
+ net2226 net951 _00335_ VPWR VGND sg13g2_mux2_1
Xhold302 _00113_ VPWR VGND net2129 sg13g2_dlygate4sd3_1
Xhold324 _00611_ VPWR VGND net2151 sg13g2_dlygate4sd3_1
Xhold335 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[6\]
+ VPWR VGND net2162 sg13g2_dlygate4sd3_1
Xhold313 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r VPWR VGND net2140
+ sg13g2_dlygate4sd3_1
X_05124_ _01854_ _01777_ i_exotiny._0013_\[2\] _01761_ i_exotiny._0015_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold357 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[18\]
+ VPWR VGND net2184 sg13g2_dlygate4sd3_1
Xhold368 _01184_ VPWR VGND net2195 sg13g2_dlygate4sd3_1
Xhold346 _01193_ VPWR VGND net2173 sg13g2_dlygate4sd3_1
X_05055_ net1221 _01753_ _01759_ _01787_ VPWR VGND sg13g2_nor3_2
XFILLER_104_439 VPWR VGND sg13g2_decap_8
Xhold379 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[15\]
+ VPWR VGND net2206 sg13g2_dlygate4sd3_1
X_08814_ net1594 VGND VPWR _00872_ i_exotiny.i_wb_spi.state_r\[13\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
Xhold1024 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[15\]
+ VPWR VGND net2851 sg13g2_dlygate4sd3_1
Xhold1013 i_exotiny._0042_\[1\] VPWR VGND net2840 sg13g2_dlygate4sd3_1
Xhold1002 _00900_ VPWR VGND net2829 sg13g2_dlygate4sd3_1
X_08745_ net1663 VGND VPWR net2549 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[8\]
+ clknet_leaf_81_clk_regs sg13g2_dfrbpq_1
Xhold1057 _00125_ VPWR VGND net2884 sg13g2_dlygate4sd3_1
Xhold1046 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[17\]
+ VPWR VGND net2873 sg13g2_dlygate4sd3_1
X_08917__1065 VPWR VGND net1485 sg13g2_tiehi
Xhold1035 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[22\]
+ VPWR VGND net2862 sg13g2_dlygate4sd3_1
X_05957_ net2406 net2729 net967 _00166_ VPWR VGND sg13g2_mux2_1
Xhold1068 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[7\]
+ VPWR VGND net2895 sg13g2_dlygate4sd3_1
Xhold1079 _00522_ VPWR VGND net2906 sg13g2_dlygate4sd3_1
XFILLER_38_261 VPWR VGND sg13g2_fill_1
X_05888_ _02473_ net2091 net1053 _00111_ VPWR VGND sg13g2_mux2_1
XFILLER_54_732 VPWR VGND sg13g2_fill_2
X_08676_ net1732 VGND VPWR _00734_ i_exotiny._0034_\[3\] clknet_leaf_122_clk_regs
+ sg13g2_dfrbpq_2
X_04908_ _01640_ i_exotiny._0077_\[2\] i_exotiny._0077_\[3\] VPWR VGND sg13g2_nand2_2
X_04839_ _01579_ _01570_ _01578_ VPWR VGND sg13g2_nand2_1
X_07627_ i_exotiny._0024_\[0\] net3105 net899 _01135_ VPWR VGND sg13g2_mux2_1
X_07558_ _03134_ VPWR _03144_ VGND net1970 _03142_ sg13g2_o21ai_1
X_06509_ _02420_ _02485_ _02620_ VPWR VGND sg13g2_nor2_2
X_07489_ VGND VPWR _01391_ net903 _01074_ _03111_ sg13g2_a21oi_1
X_09228_ net751 VGND VPWR _01283_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[18\]
+ clknet_leaf_135_clk_regs sg13g2_dfrbpq_1
X_09069__913 VPWR VGND net1333 sg13g2_tiehi
X_09159_ net823 VGND VPWR net2569 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[15\]
+ clknet_leaf_173_clk_regs sg13g2_dfrbpq_1
Xclkbuf_5_26__f_clk_regs clknet_4_13_0_clk_regs clknet_5_26__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08006__689 VPWR VGND net689 sg13g2_tiehi
X_09247__560 VPWR VGND net560 sg13g2_tiehi
XFILLER_104_951 VPWR VGND sg13g2_decap_8
Xhold891 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[30\]
+ VPWR VGND net2718 sg13g2_dlygate4sd3_1
Xhold880 _01146_ VPWR VGND net2707 sg13g2_dlygate4sd3_1
XFILLER_95_109 VPWR VGND sg13g2_fill_2
X_08568__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_103_472 VPWR VGND sg13g2_decap_8
XFILLER_89_695 VPWR VGND sg13g2_fill_1
XFILLER_76_334 VPWR VGND sg13g2_fill_2
XFILLER_92_805 VPWR VGND sg13g2_fill_1
XFILLER_67_98 VPWR VGND sg13g2_fill_2
XFILLER_91_304 VPWR VGND sg13g2_fill_1
Xhold1580 i_exotiny._0314_\[6\] VPWR VGND net3407 sg13g2_dlygate4sd3_1
X_09076__906 VPWR VGND net1326 sg13g2_tiehi
Xhold1591 _00176_ VPWR VGND net3418 sg13g2_dlygate4sd3_1
XFILLER_44_253 VPWR VGND sg13g2_fill_2
XFILLER_72_584 VPWR VGND sg13g2_fill_2
X_09254__553 VPWR VGND net553 sg13g2_tiehi
XFILLER_41_993 VPWR VGND sg13g2_fill_2
X_08306__372 VPWR VGND net372 sg13g2_tiehi
XFILLER_5_861 VPWR VGND sg13g2_decap_8
XFILLER_99_437 VPWR VGND sg13g2_decap_8
XFILLER_4_382 VPWR VGND sg13g2_fill_2
X_06860_ VGND VPWR i_exotiny._1619_\[2\] net1134 _02871_ _02870_ sg13g2_a21oi_1
Xclkbuf_leaf_184_clk_regs clknet_5_0__leaf_clk_regs clknet_leaf_184_clk_regs VPWR
+ VGND sg13g2_buf_8
X_05811_ net2214 i_exotiny._0018_\[3\] net1056 _00083_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_113_clk_regs clknet_5_25__leaf_clk_regs clknet_leaf_113_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08313__365 VPWR VGND net365 sg13g2_tiehi
X_06791_ net1133 _02811_ _02812_ _02813_ VPWR VGND sg13g2_nor3_1
X_05742_ _02378_ net3703 net1073 _00060_ VPWR VGND sg13g2_mux2_1
X_08530_ net150 VGND VPWR _00604_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[18\]
+ clknet_leaf_184_clk_regs sg13g2_dfrbpq_1
XFILLER_36_732 VPWR VGND sg13g2_fill_1
XFILLER_91_871 VPWR VGND sg13g2_fill_2
X_05673_ VGND VPWR i_exotiny._1617_\[2\] net1121 _02326_ _02325_ sg13g2_a21oi_1
XFILLER_24_927 VPWR VGND sg13g2_fill_2
X_08461_ net219 VGND VPWR net2382 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[13\]
+ clknet_leaf_163_clk_regs sg13g2_dfrbpq_1
X_04624_ _01386_ net3822 VPWR VGND sg13g2_inv_2
X_07412_ net2020 net1215 _03061_ VPWR VGND sg13g2_nor2_1
X_08392_ net286 VGND VPWR net2354 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[30\]
+ clknet_leaf_140_clk_regs sg13g2_dfrbpq_1
X_08608__1368 VPWR VGND net1788 sg13g2_tiehi
X_07343_ net3739 net1078 _03007_ VPWR VGND sg13g2_nor2_1
X_07274_ net1158 VPWR _02979_ VGND _02423_ _02978_ sg13g2_o21ai_1
X_08320__358 VPWR VGND net358 sg13g2_tiehi
X_06225_ _02544_ net2671 net945 _00377_ VPWR VGND sg13g2_mux2_1
X_09013_ net1389 VGND VPWR _01071_ i_exotiny._0327_\[1\] clknet_leaf_9_clk_regs sg13g2_dfrbpq_1
Xhold110 i_exotiny.i_wb_spi.dat_rx_r\[18\] VPWR VGND net1937 sg13g2_dlygate4sd3_1
XFILLER_3_809 VPWR VGND sg13g2_decap_8
Xhold143 i_exotiny.i_rstctl.cnt\[6\] VPWR VGND net1970 sg13g2_dlygate4sd3_1
X_06156_ net3127 net3191 net954 _00318_ VPWR VGND sg13g2_mux2_1
Xhold121 _00044_ VPWR VGND net1948 sg13g2_dlygate4sd3_1
Xhold132 i_exotiny._1924_\[31\] VPWR VGND net1959 sg13g2_dlygate4sd3_1
XFILLER_2_308 VPWR VGND sg13g2_fill_1
XFILLER_105_748 VPWR VGND sg13g2_decap_8
XFILLER_104_236 VPWR VGND sg13g2_decap_8
Xhold154 _00209_ VPWR VGND net1981 sg13g2_dlygate4sd3_1
Xhold165 _02389_ VPWR VGND net1992 sg13g2_dlygate4sd3_1
X_06087_ net2148 net3316 net955 _00263_ VPWR VGND sg13g2_mux2_1
Xhold176 _00657_ VPWR VGND net2003 sg13g2_dlygate4sd3_1
X_05107_ _01837_ _01834_ _01835_ VPWR VGND sg13g2_nand2_1
XFILLER_99_982 VPWR VGND sg13g2_decap_8
Xhold198 _01101_ VPWR VGND net2025 sg13g2_dlygate4sd3_1
X_05038_ net1221 _01757_ _01762_ _01770_ VPWR VGND sg13g2_nor3_2
Xhold187 i_exotiny._0369_\[0\] VPWR VGND net2014 sg13g2_dlygate4sd3_1
XFILLER_98_481 VPWR VGND sg13g2_decap_8
XFILLER_101_976 VPWR VGND sg13g2_decap_8
XFILLER_86_654 VPWR VGND sg13g2_fill_1
XFILLER_100_486 VPWR VGND sg13g2_decap_8
X_06989_ net2742 _02925_ net1018 _00760_ VPWR VGND sg13g2_mux2_1
XFILLER_2_1013 VPWR VGND sg13g2_decap_8
XFILLER_37_57 VPWR VGND sg13g2_fill_2
X_08728_ net1680 VGND VPWR net3184 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[23\]
+ clknet_leaf_118_clk_regs sg13g2_dfrbpq_1
X_08659_ net1738 VGND VPWR _00727_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[28\]
+ clknet_leaf_146_clk_regs sg13g2_dfrbpq_1
XFILLER_42_735 VPWR VGND sg13g2_fill_1
X_08012__682 VPWR VGND net682 sg13g2_tiehi
XFILLER_2_831 VPWR VGND sg13g2_decap_8
XFILLER_97_919 VPWR VGND sg13g2_decap_8
XFILLER_94_41 VPWR VGND sg13g2_fill_1
XFILLER_37_518 VPWR VGND sg13g2_fill_1
XFILLER_64_337 VPWR VGND sg13g2_fill_1
XFILLER_45_551 VPWR VGND sg13g2_fill_2
X_06010_ _00015_ net1105 _02499_ VPWR VGND sg13g2_nor2_1
X_07961_ net1176 VGND VPWR net3667 i_exotiny.i_wdg_top.o_wb_dat\[2\] clknet_leaf_37_clk_regs
+ sg13g2_dfrbpq_2
X_06912_ net3466 i_exotiny.core_res_en_n _02911_ _02912_ VPWR VGND sg13g2_a21o_1
XFILLER_96_963 VPWR VGND sg13g2_decap_8
X_07892_ i_exotiny._0021_\[1\] net881 _03228_ _03231_ VPWR VGND sg13g2_mux2_1
XFILLER_83_624 VPWR VGND sg13g2_fill_2
X_06843_ net3680 net1097 _02857_ VPWR VGND sg13g2_nor2_1
XFILLER_67_153 VPWR VGND sg13g2_fill_1
XFILLER_83_657 VPWR VGND sg13g2_fill_2
X_06774_ net2042 net1100 _02799_ VPWR VGND sg13g2_nor2_1
X_05725_ net1928 net1058 _02365_ VPWR VGND sg13g2_nor2_1
X_09059__923 VPWR VGND net1343 sg13g2_tiehi
X_08513_ net167 VGND VPWR net2286 i_exotiny._0043_\[1\] clknet_leaf_177_clk_regs sg13g2_dfrbpq_2
Xclkbuf_4_10_0_clk_regs clknet_0_clk_regs clknet_4_10_0_clk_regs VPWR VGND sg13g2_buf_8
Xclkbuf_leaf_81_clk_regs clknet_5_27__leaf_clk_regs clknet_leaf_81_clk_regs VPWR VGND
+ sg13g2_buf_8
X_05656_ net1122 net1939 _02313_ VPWR VGND sg13g2_nor2b_1
X_08444_ net238 VGND VPWR _00518_ i_exotiny._2025_\[6\] clknet_leaf_28_clk_regs sg13g2_dfrbpq_2
XFILLER_51_554 VPWR VGND sg13g2_fill_1
XFILLER_11_418 VPWR VGND sg13g2_fill_2
X_08375_ net303 VGND VPWR net2651 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[13\]
+ clknet_leaf_138_clk_regs sg13g2_dfrbpq_1
X_04607_ VPWR _01369_ net2037 VGND sg13g2_inv_1
XFILLER_23_26 VPWR VGND sg13g2_fill_2
X_05587_ _02261_ _02258_ _02262_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_10_clk_regs clknet_5_3__leaf_clk_regs clknet_leaf_10_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07326_ net1214 _02988_ _02990_ VPWR VGND sg13g2_nor2_1
X_09268__91 VPWR VGND net91 sg13g2_tiehi
X_07257_ net2759 net2309 net1004 _00980_ VPWR VGND sg13g2_mux2_1
XFILLER_105_501 VPWR VGND sg13g2_decap_8
X_06208_ net2375 net2863 net947 _00363_ VPWR VGND sg13g2_mux2_1
X_07188_ VGND VPWR _01366_ _02956_ _00926_ net3742 sg13g2_a21oi_1
X_09066__916 VPWR VGND net1336 sg13g2_tiehi
XFILLER_3_7 VPWR VGND sg13g2_decap_8
X_06139_ net2664 net3011 net1045 _00308_ VPWR VGND sg13g2_mux2_1
XFILLER_105_578 VPWR VGND sg13g2_decap_8
X_09244__563 VPWR VGND net563 sg13g2_tiehi
XFILLER_87_985 VPWR VGND sg13g2_decap_8
XFILLER_100_283 VPWR VGND sg13g2_decap_8
XFILLER_104_84 VPWR VGND sg13g2_fill_1
X_08654__1323 VPWR VGND net1743 sg13g2_tiehi
X_09073__909 VPWR VGND net1329 sg13g2_tiehi
XFILLER_55_882 VPWR VGND sg13g2_fill_1
X_09251__556 VPWR VGND net556 sg13g2_tiehi
XFILLER_11_974 VPWR VGND sg13g2_decap_8
XFILLER_7_912 VPWR VGND sg13g2_decap_8
X_08303__375 VPWR VGND net375 sg13g2_tiehi
XFILLER_7_989 VPWR VGND sg13g2_decap_8
X_08876__1106 VPWR VGND net1526 sg13g2_tiehi
X_08912__1070 VPWR VGND net1490 sg13g2_tiehi
XFILLER_2_650 VPWR VGND sg13g2_fill_1
XFILLER_96_204 VPWR VGND sg13g2_fill_1
XFILLER_36_7 VPWR VGND sg13g2_decap_8
X_07958__698 VPWR VGND net698 sg13g2_tiehi
XFILLER_92_410 VPWR VGND sg13g2_fill_1
XFILLER_49_164 VPWR VGND sg13g2_fill_2
XFILLER_93_977 VPWR VGND sg13g2_decap_8
X_08310__368 VPWR VGND net368 sg13g2_tiehi
XFILLER_92_476 VPWR VGND sg13g2_fill_2
XFILLER_18_584 VPWR VGND sg13g2_fill_1
X_06490_ net3101 net2876 net1025 _00571_ VPWR VGND sg13g2_mux2_1
X_05510_ _02200_ VPWR i_exotiny._1611_\[17\] VGND net1074 _02202_ sg13g2_o21ai_1
X_05441_ _02150_ _02149_ i_exotiny._1617_\[0\] _02148_ i_exotiny._1612_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_08160_ net518 VGND VPWR _00241_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[24\]
+ clknet_leaf_120_clk_regs sg13g2_dfrbpq_1
X_07111_ net1288 net1861 _00861_ VPWR VGND sg13g2_and2_1
X_05372_ VGND VPWR _02092_ _02093_ _02094_ _02075_ sg13g2_a21oi_1
XFILLER_20_259 VPWR VGND sg13g2_fill_2
X_08091_ net603 VGND VPWR net2813 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[28\]
+ clknet_leaf_86_clk_regs sg13g2_dfrbpq_1
X_07042_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[12\]
+ net2548 net1013 _00803_ VPWR VGND sg13g2_mux2_1
Xclkload30 clkload30/Y clknet_leaf_51_clk_regs VPWR VGND sg13g2_inv_2
Xclkload41 VPWR clkload41/Y clknet_leaf_106_clk_regs VGND sg13g2_inv_1
XFILLER_102_504 VPWR VGND sg13g2_decap_8
X_08993_ net1409 VGND VPWR net2041 i_exotiny._1160_\[14\] clknet_leaf_162_clk_regs
+ sg13g2_dfrbpq_1
X_08732__1256 VPWR VGND net1676 sg13g2_tiehi
X_07944_ net88 VGND VPWR net3755 i_exotiny._1660_ clknet_leaf_27_clk_regs sg13g2_dfrbpq_2
XFILLER_56_624 VPWR VGND sg13g2_fill_1
X_07875_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[13\]
+ net2211 net978 _01342_ VPWR VGND sg13g2_mux2_1
X_06826_ VGND VPWR net1099 _02841_ _00680_ _02842_ sg13g2_a21oi_1
XFILLER_93_1012 VPWR VGND sg13g2_decap_8
X_06757_ VGND VPWR _01412_ net1191 _02784_ _02783_ sg13g2_a21oi_1
X_05708_ net1115 i_exotiny._1924_\[27\] _02352_ VPWR VGND sg13g2_nor2b_1
X_06688_ _02593_ _02722_ _02723_ _02725_ VPWR VGND sg13g2_nor3_1
XFILLER_24_543 VPWR VGND sg13g2_fill_2
X_08954__1028 VPWR VGND net1448 sg13g2_tiehi
X_05639_ net1909 net1065 _02300_ VPWR VGND sg13g2_nor2_1
X_08427_ net258 VGND VPWR _00501_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[26\]
+ clknet_leaf_96_clk_regs sg13g2_dfrbpq_1
XFILLER_24_565 VPWR VGND sg13g2_fill_1
Xclkload2 clkload2/Y clknet_5_11__leaf_clk_regs VPWR VGND sg13g2_inv_2
X_08358_ net320 VGND VPWR net2384 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[28\]
+ clknet_leaf_95_clk_regs sg13g2_dfrbpq_1
X_07309_ net872 net3013 _02978_ _02983_ VPWR VGND sg13g2_mux2_1
X_08289_ net389 VGND VPWR _00370_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[23\]
+ clknet_leaf_100_clk_regs sg13g2_dfrbpq_1
XFILLER_4_904 VPWR VGND sg13g2_decap_8
XFILLER_106_832 VPWR VGND sg13g2_decap_8
XFILLER_59_33 VPWR VGND sg13g2_fill_1
XFILLER_105_375 VPWR VGND sg13g2_decap_8
Xfanout1204 net1206 net1204 VPWR VGND sg13g2_buf_8
Xfanout1226 net1227 net1226 VPWR VGND sg13g2_buf_8
Xfanout1215 net1217 net1215 VPWR VGND sg13g2_buf_8
X_08708__1280 VPWR VGND net1700 sg13g2_tiehi
Xfanout1237 i_exotiny._0079_\[4\] net1237 VPWR VGND sg13g2_buf_8
Xfanout1248 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[5\]
+ net1248 VPWR VGND sg13g2_buf_8
X_08118__576 VPWR VGND net576 sg13g2_tiehi
Xfanout1259 net3812 net1259 VPWR VGND sg13g2_buf_2
XFILLER_75_955 VPWR VGND sg13g2_fill_1
XFILLER_19_337 VPWR VGND sg13g2_fill_1
XFILLER_62_616 VPWR VGND sg13g2_fill_1
XFILLER_47_668 VPWR VGND sg13g2_decap_4
XFILLER_90_947 VPWR VGND sg13g2_decap_8
XFILLER_74_487 VPWR VGND sg13g2_fill_1
X_08603__1373 VPWR VGND net1793 sg13g2_tiehi
XFILLER_43_863 VPWR VGND sg13g2_fill_2
XFILLER_15_565 VPWR VGND sg13g2_fill_1
X_08810__1178 VPWR VGND net1598 sg13g2_tiehi
X_08125__569 VPWR VGND net569 sg13g2_tiehi
Xhold709 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[27\]
+ VPWR VGND net2536 sg13g2_dlygate4sd3_1
XFILLER_40_90 VPWR VGND sg13g2_fill_1
XFILLER_97_502 VPWR VGND sg13g2_decap_8
XFILLER_3_970 VPWR VGND sg13g2_decap_8
XFILLER_34_4 VPWR VGND sg13g2_decap_8
XFILLER_69_248 VPWR VGND sg13g2_fill_2
X_05990_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[16\]
+ net2343 net1050 _00192_ VPWR VGND sg13g2_mux2_1
Xhold1409 _03174_ VPWR VGND net3236 sg13g2_dlygate4sd3_1
X_04941_ _01659_ _01662_ _01672_ _01673_ VPWR VGND sg13g2_nor3_2
XFILLER_65_443 VPWR VGND sg13g2_fill_2
X_07660_ net2296 _03191_ net896 _01165_ VPWR VGND sg13g2_mux2_1
X_04872_ net1250 _01427_ net1248 _01604_ VPWR VGND sg13g2_nand3_1
XFILLER_92_284 VPWR VGND sg13g2_decap_8
X_07591_ net1206 net2029 _03165_ _01122_ VPWR VGND sg13g2_nor3_1
X_06611_ net3358 net1152 _02664_ VPWR VGND sg13g2_nor2_1
X_09056__926 VPWR VGND net1346 sg13g2_tiehi
X_06542_ net2150 _02623_ net929 _00615_ VPWR VGND sg13g2_mux2_1
XFILLER_61_671 VPWR VGND sg13g2_fill_1
X_09261_ net239 VGND VPWR net3421 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[19\]
+ clknet_leaf_129_clk_regs sg13g2_dfrbpq_1
XFILLER_33_351 VPWR VGND sg13g2_fill_1
X_06473_ net3351 net2703 net1024 _00554_ VPWR VGND sg13g2_mux2_1
X_08212_ net465 VGND VPWR net2603 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[11\]
+ clknet_leaf_150_clk_regs sg13g2_dfrbpq_1
X_09192_ net789 VGND VPWR net2582 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[14\]
+ clknet_leaf_79_clk_regs sg13g2_dfrbpq_1
X_05424_ _02133_ net1230 _02131_ VPWR VGND sg13g2_xnor2_1
X_05355_ _02077_ _01400_ _01375_ i_exotiny._2034_\[1\] _00015_ VPWR VGND sg13g2_a22oi_1
X_08143_ net542 VGND VPWR _00224_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[7\]
+ clknet_leaf_118_clk_regs sg13g2_dfrbpq_1
X_08074_ net620 VGND VPWR net2823 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[11\]
+ clknet_leaf_93_clk_regs sg13g2_dfrbpq_1
XFILLER_106_139 VPWR VGND sg13g2_decap_8
X_05286_ VGND VPWR _01750_ _02011_ _02012_ net1108 sg13g2_a21oi_1
X_07025_ net2083 _02930_ net918 _00791_ VPWR VGND sg13g2_mux2_1
X_09263__235 VPWR VGND net235 sg13g2_tiehi
XFILLER_102_301 VPWR VGND sg13g2_decap_8
X_09063__919 VPWR VGND net1339 sg13g2_tiehi
XFILLER_1_929 VPWR VGND sg13g2_decap_8
XFILLER_103_846 VPWR VGND sg13g2_decap_8
Xhold14 i_exotiny.i_wb_spi.state_r\[15\] VPWR VGND net1841 sg13g2_dlygate4sd3_1
XFILLER_102_378 VPWR VGND sg13g2_decap_8
Xhold25 i_exotiny.i_wb_spi.state_r\[20\] VPWR VGND net1852 sg13g2_dlygate4sd3_1
Xhold36 i_exotiny.i_wb_spi.state_r\[1\] VPWR VGND net1863 sg13g2_dlygate4sd3_1
Xhold47 _00079_ VPWR VGND net1874 sg13g2_dlygate4sd3_1
X_09241__566 VPWR VGND net566 sg13g2_tiehi
Xhold1910 i_exotiny._0369_\[18\] VPWR VGND net3737 sg13g2_dlygate4sd3_1
X_08976_ net1426 VGND VPWR _01034_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[1\]
+ clknet_leaf_15_clk_regs sg13g2_dfrbpq_2
Xhold58 i_exotiny.i_wdg_top.clk_div_inst.cnt\[3\] VPWR VGND net1885 sg13g2_dlygate4sd3_1
Xhold1954 _02072_ VPWR VGND net3781 sg13g2_dlygate4sd3_1
Xhold69 _00032_ VPWR VGND net1896 sg13g2_dlygate4sd3_1
X_07927_ net721 VGND VPWR net1958 i_exotiny._1924_\[20\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
XFILLER_57_944 VPWR VGND sg13g2_fill_2
Xhold1921 _00691_ VPWR VGND net3748 sg13g2_dlygate4sd3_1
Xhold1932 i_exotiny._0369_\[12\] VPWR VGND net3759 sg13g2_dlygate4sd3_1
Xhold1943 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[1\]
+ VPWR VGND net3770 sg13g2_dlygate4sd3_1
Xhold1965 _02409_ VPWR VGND net3792 sg13g2_dlygate4sd3_1
Xhold1987 i_exotiny.i_wb_spi.cnt_presc_r\[2\] VPWR VGND net3814 sg13g2_dlygate4sd3_1
XFILLER_57_977 VPWR VGND sg13g2_fill_1
X_07858_ net2592 net875 _03222_ _03227_ VPWR VGND sg13g2_mux2_1
Xhold1976 _03020_ VPWR VGND net3803 sg13g2_dlygate4sd3_1
X_06809_ i_exotiny._0369_\[18\] net1188 _02828_ VPWR VGND sg13g2_nor2_1
X_07789_ net3249 net3508 net892 _01268_ VPWR VGND sg13g2_mux2_1
XFILLER_28_167 VPWR VGND sg13g2_fill_1
Xhold1998 i_exotiny._0079_\[3\] VPWR VGND net3825 sg13g2_dlygate4sd3_1
XFILLER_37_690 VPWR VGND sg13g2_fill_2
XFILLER_40_844 VPWR VGND sg13g2_fill_1
X_08300__378 VPWR VGND net378 sg13g2_tiehi
XFILLER_4_778 VPWR VGND sg13g2_decap_8
XFILLER_105_172 VPWR VGND sg13g2_decap_8
Xfanout1012 _02948_ net1012 VPWR VGND sg13g2_buf_8
Xfanout1001 net1002 net1001 VPWR VGND sg13g2_buf_8
Xfanout1056 _02424_ net1056 VPWR VGND sg13g2_buf_8
Xfanout1023 net1024 net1023 VPWR VGND sg13g2_buf_8
XFILLER_0_973 VPWR VGND sg13g2_decap_8
Xfanout1034 net1037 net1034 VPWR VGND sg13g2_buf_8
Xfanout1045 _02527_ net1045 VPWR VGND sg13g2_buf_8
Xfanout1089 net1090 net1089 VPWR VGND sg13g2_buf_1
Xfanout1067 _02273_ net1067 VPWR VGND sg13g2_buf_8
Xfanout1078 _02991_ net1078 VPWR VGND sg13g2_buf_8
XFILLER_19_134 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_138_clk_regs clknet_5_17__leaf_clk_regs clknet_leaf_138_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_16_896 VPWR VGND sg13g2_fill_2
XFILLER_30_387 VPWR VGND sg13g2_fill_1
X_05140_ VGND VPWR _01750_ _01869_ _01870_ net1108 sg13g2_a21oi_1
Xhold517 _00192_ VPWR VGND net2344 sg13g2_dlygate4sd3_1
Xhold506 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[27\]
+ VPWR VGND net2333 sg13g2_dlygate4sd3_1
XFILLER_7_572 VPWR VGND sg13g2_fill_2
XFILLER_7_561 VPWR VGND sg13g2_fill_1
XFILLER_83_1000 VPWR VGND sg13g2_decap_8
X_08199__478 VPWR VGND net478 sg13g2_tiehi
Xhold528 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[28\]
+ VPWR VGND net2355 sg13g2_dlygate4sd3_1
Xhold539 _01334_ VPWR VGND net2366 sg13g2_dlygate4sd3_1
X_05071_ _01803_ _01787_ i_exotiny._0031_\[3\] _01776_ i_exotiny._0021_\[3\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_97_310 VPWR VGND sg13g2_decap_8
X_08830_ net1578 VGND VPWR _00888_ i_exotiny.i_wb_spi.state_r\[29\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_100_805 VPWR VGND sg13g2_decap_8
XFILLER_98_888 VPWR VGND sg13g2_decap_8
Xhold1206 _00715_ VPWR VGND net3033 sg13g2_dlygate4sd3_1
XFILLER_25_0 VPWR VGND sg13g2_fill_2
XFILLER_97_387 VPWR VGND sg13g2_decap_8
X_08761_ net1647 VGND VPWR _00819_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[24\]
+ clknet_leaf_80_clk_regs sg13g2_dfrbpq_1
X_05973_ _02493_ net1139 net1167 _02494_ VPWR VGND sg13g2_a21o_1
Xhold1239 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[30\]
+ VPWR VGND net3066 sg13g2_dlygate4sd3_1
Xhold1228 _00603_ VPWR VGND net3055 sg13g2_dlygate4sd3_1
Xhold1217 i_exotiny._0014_\[3\] VPWR VGND net3044 sg13g2_dlygate4sd3_1
X_08692_ net1716 VGND VPWR _00750_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[19\]
+ clknet_leaf_105_clk_regs sg13g2_dfrbpq_1
X_07712_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[13\]
+ net2545 net997 _01208_ VPWR VGND sg13g2_mux2_1
X_04924_ _01656_ _01648_ i_exotiny._0033_\[3\] _01646_ i_exotiny._0017_\[3\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_93_582 VPWR VGND sg13g2_fill_2
X_04855_ VGND VPWR net3618 _01570_ _01591_ net1072 sg13g2_a21oi_1
XFILLER_65_251 VPWR VGND sg13g2_fill_2
X_07643_ net2785 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[20\]
+ net899 _01151_ VPWR VGND sg13g2_mux2_1
X_07574_ net1204 _03153_ _03154_ _01116_ VPWR VGND sg13g2_nor3_1
XFILLER_81_788 VPWR VGND sg13g2_fill_2
X_04786_ net1273 _01437_ _01536_ VPWR VGND sg13g2_nor2_1
X_06525_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[14\]
+ net2184 net929 _00600_ VPWR VGND sg13g2_mux2_1
XFILLER_34_682 VPWR VGND sg13g2_fill_1
X_08871__1111 VPWR VGND net1531 sg13g2_tiehi
X_06456_ net3172 net2955 net934 _00543_ VPWR VGND sg13g2_mux2_1
X_09244_ net563 VGND VPWR net2163 i_exotiny._0022_\[2\] clknet_leaf_123_clk_regs sg13g2_dfrbpq_2
X_05407_ net1113 _02118_ _02119_ i_exotiny._2043_\[6\] VPWR VGND sg13g2_nor3_1
X_09175_ net807 VGND VPWR _01230_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[31\]
+ clknet_leaf_173_clk_regs sg13g2_dfrbpq_1
X_08108__586 VPWR VGND net586 sg13g2_tiehi
X_06387_ net1225 net3648 _00508_ VPWR VGND sg13g2_nor2_1
X_08126_ net568 VGND VPWR _00207_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[31\]
+ clknet_leaf_123_clk_regs sg13g2_dfrbpq_1
Xclkbuf_5_25__f_clk_regs clknet_4_12_0_clk_regs clknet_5_25__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_05338_ i_exotiny._1266_ VPWR _02062_ VGND _01459_ _01678_ sg13g2_o21ai_1
X_08057_ net637 VGND VPWR _00138_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[26\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
X_05269_ _01995_ _01776_ i_exotiny._0021_\[0\] _01760_ i_exotiny._0014_\[0\] VPWR
+ VGND sg13g2_a22oi_1
Xoutput37 net37 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_726 VPWR VGND sg13g2_decap_8
Xoutput26 net26 uio_out[0] VPWR VGND sg13g2_buf_1
X_07008_ net2872 net2645 net922 _00775_ VPWR VGND sg13g2_mux2_1
XFILLER_89_877 VPWR VGND sg13g2_fill_1
XFILLER_102_175 VPWR VGND sg13g2_decap_8
X_09178__803 VPWR VGND net803 sg13g2_tiehi
X_08959_ net1443 VGND VPWR _01017_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[25\]
+ clknet_leaf_60_clk_regs sg13g2_dfrbpq_1
XFILLER_5_1022 VPWR VGND sg13g2_decap_8
Xhold1751 i_exotiny.i_wdg_top.clk_div_inst.cnt\[11\] VPWR VGND net3578 sg13g2_dlygate4sd3_1
Xhold1740 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data[0]
+ VPWR VGND net3567 sg13g2_dlygate4sd3_1
Xhold1762 i_exotiny.i_wb_spi.dat_rx_r\[0\] VPWR VGND net3589 sg13g2_dlygate4sd3_1
Xhold1795 i_exotiny._1615_\[2\] VPWR VGND net3622 sg13g2_dlygate4sd3_1
Xhold1773 i_exotiny.i_wb_spi.dat_rx_r\[21\] VPWR VGND net3600 sg13g2_dlygate4sd3_1
XFILLER_57_785 VPWR VGND sg13g2_fill_1
X_08115__579 VPWR VGND net579 sg13g2_tiehi
Xhold1784 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data[0]
+ VPWR VGND net3611 sg13g2_dlygate4sd3_1
X_09039__943 VPWR VGND net1363 sg13g2_tiehi
XFILLER_72_77 VPWR VGND sg13g2_fill_1
XFILLER_71_287 VPWR VGND sg13g2_fill_1
XFILLER_9_804 VPWR VGND sg13g2_fill_2
X_09046__936 VPWR VGND net1356 sg13g2_tiehi
XFILLER_39_207 VPWR VGND sg13g2_fill_1
XFILLER_67_538 VPWR VGND sg13g2_fill_2
XFILLER_67_527 VPWR VGND sg13g2_fill_1
XFILLER_0_770 VPWR VGND sg13g2_decap_8
X_09043__1150 VPWR VGND net1570 sg13g2_tiehi
XFILLER_36_936 VPWR VGND sg13g2_fill_1
XFILLER_47_295 VPWR VGND sg13g2_fill_1
X_04640_ _01402_ net3780 VPWR VGND sg13g2_inv_2
X_09053__929 VPWR VGND net1349 sg13g2_tiehi
X_07290_ net2954 net2846 net911 _01007_ VPWR VGND sg13g2_mux2_1
X_06310_ net2426 net3429 net1035 _00447_ VPWR VGND sg13g2_mux2_1
X_06241_ net2914 net2415 net1039 _00390_ VPWR VGND sg13g2_mux2_1
X_06172_ net2109 net2554 net953 _00334_ VPWR VGND sg13g2_mux2_1
XFILLER_11_1027 VPWR VGND sg13g2_fill_2
XFILLER_11_1016 VPWR VGND sg13g2_decap_8
Xhold325 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[16\]
+ VPWR VGND net2152 sg13g2_dlygate4sd3_1
Xhold303 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[22\]
+ VPWR VGND net2130 sg13g2_dlygate4sd3_1
Xhold314 _00249_ VPWR VGND net2141 sg13g2_dlygate4sd3_1
X_05123_ _01853_ _01789_ i_exotiny._0024_\[2\] _01765_ i_exotiny._0027_\[2\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_104_418 VPWR VGND sg13g2_decap_8
XFILLER_89_107 VPWR VGND sg13g2_fill_1
Xhold369 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[26\]
+ VPWR VGND net2196 sg13g2_dlygate4sd3_1
Xhold347 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[4\]
+ VPWR VGND net2174 sg13g2_dlygate4sd3_1
Xhold358 _00600_ VPWR VGND net2185 sg13g2_dlygate4sd3_1
Xhold336 _01299_ VPWR VGND net2163 sg13g2_dlygate4sd3_1
X_05054_ net1236 _01754_ _01756_ _01786_ VPWR VGND sg13g2_nor3_2
Xclkbuf_leaf_35_clk_regs clknet_5_9__leaf_clk_regs clknet_leaf_35_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_98_685 VPWR VGND sg13g2_fill_1
XFILLER_98_674 VPWR VGND sg13g2_fill_1
Xhold1003 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[24\]
+ VPWR VGND net2830 sg13g2_dlygate4sd3_1
X_08813_ net1595 VGND VPWR net1850 i_exotiny.i_wb_spi.state_r\[12\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
Xhold1014 i_exotiny._0315_\[24\] VPWR VGND net2841 sg13g2_dlygate4sd3_1
X_08744_ net1664 VGND VPWR net3110 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[7\]
+ clknet_leaf_81_clk_regs sg13g2_dfrbpq_1
X_05956_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[21\]
+ net2458 net970 _00165_ VPWR VGND sg13g2_mux2_1
XFILLER_85_368 VPWR VGND sg13g2_fill_2
Xhold1025 _00490_ VPWR VGND net2852 sg13g2_dlygate4sd3_1
Xhold1036 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[16\]
+ VPWR VGND net2863 sg13g2_dlygate4sd3_1
Xhold1058 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[23\]
+ VPWR VGND net2885 sg13g2_dlygate4sd3_1
Xhold1047 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[16\]
+ VPWR VGND net2874 sg13g2_dlygate4sd3_1
Xhold1069 _00115_ VPWR VGND net2896 sg13g2_dlygate4sd3_1
X_04907_ _01639_ _01638_ i_exotiny._0029_\[3\] _01637_ i_exotiny._0024_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_05887_ net2639 net872 _02421_ _02473_ VPWR VGND sg13g2_mux2_1
X_08675_ net1733 VGND VPWR net2244 i_exotiny._0034_\[2\] clknet_leaf_104_clk_regs
+ sg13g2_dfrbpq_2
X_07942__86 VPWR VGND net86 sg13g2_tiehi
Xclkbuf_5_9__f_clk_regs clknet_4_4_0_clk_regs clknet_5_9__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_04838_ net1187 _01485_ _01578_ VPWR VGND sg13g2_nor2_2
X_07626_ _03187_ net1141 net1168 _03188_ VPWR VGND sg13g2_a21o_2
X_07557_ _03142_ _03143_ _01110_ VPWR VGND sg13g2_nor2_1
X_04769_ net3830 _01519_ _01520_ VPWR VGND sg13g2_and2_1
X_06508_ _02619_ net3117 net1024 _00585_ VPWR VGND sg13g2_mux2_1
XFILLER_21_151 VPWR VGND sg13g2_fill_2
X_07488_ net3670 net907 _03111_ VPWR VGND sg13g2_nor2_1
X_06439_ net2609 net2905 net937 _00526_ VPWR VGND sg13g2_mux2_1
X_09227_ net752 VGND VPWR net2626 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[17\]
+ clknet_leaf_129_clk_regs sg13g2_dfrbpq_1
X_09158_ net824 VGND VPWR net2423 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[14\]
+ clknet_leaf_148_clk_regs sg13g2_dfrbpq_1
X_08109_ net585 VGND VPWR _00190_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[14\]
+ clknet_leaf_122_clk_regs sg13g2_dfrbpq_1
X_09089_ net1313 VGND VPWR _01144_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[9\]
+ clknet_leaf_142_clk_regs sg13g2_dfrbpq_1
XFILLER_101_4 VPWR VGND sg13g2_fill_2
XFILLER_104_930 VPWR VGND sg13g2_decap_8
Xhold870 _01258_ VPWR VGND net2697 sg13g2_dlygate4sd3_1
Xhold881 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[12\]
+ VPWR VGND net2708 sg13g2_dlygate4sd3_1
XFILLER_103_451 VPWR VGND sg13g2_decap_8
XFILLER_88_151 VPWR VGND sg13g2_fill_2
Xhold892 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[27\]
+ VPWR VGND net2719 sg13g2_dlygate4sd3_1
XFILLER_88_173 VPWR VGND sg13g2_fill_2
XFILLER_77_836 VPWR VGND sg13g2_fill_2
XFILLER_1_589 VPWR VGND sg13g2_fill_1
XFILLER_67_77 VPWR VGND sg13g2_fill_2
Xhold1570 i_exotiny._0036_\[2\] VPWR VGND net3397 sg13g2_dlygate4sd3_1
X_08745__1243 VPWR VGND net1663 sg13g2_tiehi
Xhold1592 i_exotiny._0035_\[1\] VPWR VGND net3419 sg13g2_dlygate4sd3_1
Xhold1581 _00630_ VPWR VGND net3408 sg13g2_dlygate4sd3_1
XFILLER_29_284 VPWR VGND sg13g2_fill_2
X_08189__488 VPWR VGND net488 sg13g2_tiehi
XFILLER_9_623 VPWR VGND sg13g2_fill_1
XFILLER_5_840 VPWR VGND sg13g2_decap_8
X_08967__1015 VPWR VGND net1435 sg13g2_tiehi
XFILLER_99_416 VPWR VGND sg13g2_decap_8
X_05810_ net2802 net3282 net1056 _00082_ VPWR VGND sg13g2_mux2_1
X_06790_ net1171 VPWR _02812_ VGND net2432 net1185 sg13g2_o21ai_1
X_07990__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_82_338 VPWR VGND sg13g2_fill_2
X_05741_ _02375_ VPWR _02378_ VGND net1118 _02377_ sg13g2_o21ai_1
Xclkbuf_leaf_153_clk_regs clknet_5_18__leaf_clk_regs clknet_leaf_153_clk_regs VPWR
+ VGND sg13g2_buf_8
X_05672_ net1123 net1901 _02325_ VPWR VGND sg13g2_nor2b_1
X_08460_ net220 VGND VPWR _00534_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[12\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_1
XFILLER_50_213 VPWR VGND sg13g2_fill_2
X_08391_ net287 VGND VPWR net3148 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[29\]
+ clknet_leaf_139_clk_regs sg13g2_dfrbpq_1
X_07411_ net1080 net2101 _03060_ _01047_ VPWR VGND sg13g2_a21o_1
X_04623_ net1267 _01385_ VPWR VGND sg13g2_inv_4
X_07342_ VGND VPWR net3712 net1212 _03006_ _03005_ sg13g2_a21oi_1
XFILLER_31_460 VPWR VGND sg13g2_fill_1
X_07273_ _02978_ _02476_ VPWR VGND _02420_ sg13g2_nand2b_2
X_08616__1360 VPWR VGND net1780 sg13g2_tiehi
X_06224_ i_exotiny._0033_\[2\] net878 _02540_ _02544_ VPWR VGND sg13g2_mux2_1
X_09012_ net1390 VGND VPWR _01070_ i_exotiny._0327_\[0\] clknet_leaf_9_clk_regs sg13g2_dfrbpq_2
X_06155_ i_exotiny._0028_\[3\] net3102 net950 _00317_ VPWR VGND sg13g2_mux2_1
Xhold100 _00047_ VPWR VGND net1927 sg13g2_dlygate4sd3_1
XFILLER_105_727 VPWR VGND sg13g2_decap_8
Xhold144 _01111_ VPWR VGND net1971 sg13g2_dlygate4sd3_1
Xhold111 _00946_ VPWR VGND net1938 sg13g2_dlygate4sd3_1
Xhold133 _00056_ VPWR VGND net1960 sg13g2_dlygate4sd3_1
X_08105__589 VPWR VGND net589 sg13g2_tiehi
X_05106_ _01834_ _01835_ _01836_ VPWR VGND sg13g2_and2_1
Xhold122 i_exotiny._1160_\[3\] VPWR VGND net1949 sg13g2_dlygate4sd3_1
X_08823__1165 VPWR VGND net1585 sg13g2_tiehi
XFILLER_104_215 VPWR VGND sg13g2_decap_8
Xhold166 _00065_ VPWR VGND net1993 sg13g2_dlygate4sd3_1
X_08005__690 VPWR VGND net690 sg13g2_tiehi
Xhold177 i_exotiny._1924_\[16\] VPWR VGND net2004 sg13g2_dlygate4sd3_1
Xhold155 i_exotiny._1924_\[26\] VPWR VGND net1982 sg13g2_dlygate4sd3_1
X_06086_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[12\]
+ net2844 net956 _00262_ VPWR VGND sg13g2_mux2_1
XFILLER_99_961 VPWR VGND sg13g2_decap_8
X_09029__953 VPWR VGND net1373 sg13g2_tiehi
Xhold199 i_exotiny._1160_\[6\] VPWR VGND net2026 sg13g2_dlygate4sd3_1
X_05037_ _01753_ _01768_ _01769_ VPWR VGND sg13g2_nor2_2
Xhold188 _00514_ VPWR VGND net2015 sg13g2_dlygate4sd3_1
XFILLER_98_460 VPWR VGND sg13g2_decap_8
XFILLER_101_955 VPWR VGND sg13g2_decap_8
XFILLER_85_121 VPWR VGND sg13g2_fill_2
XFILLER_100_465 VPWR VGND sg13g2_decap_8
XFILLER_58_379 VPWR VGND sg13g2_fill_2
X_06988_ net3104 net883 _02922_ _02925_ VPWR VGND sg13g2_mux2_1
XFILLER_39_560 VPWR VGND sg13g2_decap_4
X_05939_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[4\]
+ net2319 net968 _00148_ VPWR VGND sg13g2_mux2_1
XFILLER_27_733 VPWR VGND sg13g2_fill_1
XFILLER_37_69 VPWR VGND sg13g2_fill_1
X_08727_ net1681 VGND VPWR net2112 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[22\]
+ clknet_leaf_121_clk_regs sg13g2_dfrbpq_1
X_08658_ net1739 VGND VPWR _00726_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[27\]
+ clknet_leaf_147_clk_regs sg13g2_dfrbpq_1
XFILLER_27_777 VPWR VGND sg13g2_fill_1
X_07609_ i_exotiny._0000_ VPWR _03177_ VGND net3722 _03175_ sg13g2_o21ai_1
XFILLER_23_950 VPWR VGND sg13g2_fill_1
X_08589_ net1807 VGND VPWR _00661_ i_exotiny._6090_\[1\] clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
X_09036__946 VPWR VGND net1366 sg13g2_tiehi
XFILLER_41_279 VPWR VGND sg13g2_fill_2
XFILLER_78_32 VPWR VGND sg13g2_fill_2
XFILLER_2_810 VPWR VGND sg13g2_decap_8
X_09082__900 VPWR VGND net1320 sg13g2_tiehi
XFILLER_77_622 VPWR VGND sg13g2_fill_1
X_07974__115 VPWR VGND net115 sg13g2_tiehi
XFILLER_2_887 VPWR VGND sg13g2_decap_8
XFILLER_49_346 VPWR VGND sg13g2_fill_1
XFILLER_73_883 VPWR VGND sg13g2_fill_1
XFILLER_72_393 VPWR VGND sg13g2_fill_2
XFILLER_17_298 VPWR VGND sg13g2_fill_2
XFILLER_9_453 VPWR VGND sg13g2_fill_2
X_07960_ net1175 VGND VPWR net3554 i_exotiny.i_wdg_top.o_wb_dat\[1\] clknet_leaf_37_clk_regs
+ sg13g2_dfrbpq_2
X_06911_ net2298 net1970 _02909_ _02910_ _02911_ VPWR VGND sg13g2_nor4_1
XFILLER_96_942 VPWR VGND sg13g2_decap_8
XFILLER_67_110 VPWR VGND sg13g2_fill_2
X_07891_ net2253 _03230_ net978 _01357_ VPWR VGND sg13g2_mux2_1
XFILLER_95_474 VPWR VGND sg13g2_fill_1
X_06842_ VGND VPWR net3620 net1132 _02856_ _02855_ sg13g2_a21oi_1
XFILLER_55_305 VPWR VGND sg13g2_fill_1
X_06773_ VGND VPWR net2063 net1135 _02798_ _02797_ sg13g2_a21oi_1
X_05724_ VGND VPWR i_exotiny._1618_\[3\] net1115 _02364_ _02363_ sg13g2_a21oi_1
X_08512_ net168 VGND VPWR _00586_ i_exotiny._0043_\[0\] clknet_leaf_175_clk_regs sg13g2_dfrbpq_2
X_08570__64 VPWR VGND net64 sg13g2_tiehi
X_05655_ net1963 net1063 _02312_ VPWR VGND sg13g2_nor2_1
X_08443_ net240 VGND VPWR _00517_ i_exotiny._2025_\[5\] clknet_leaf_29_clk_regs sg13g2_dfrbpq_2
X_04606_ VPWR _01368_ net3466 VGND sg13g2_inv_1
X_08374_ net304 VGND VPWR net2326 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[12\]
+ clknet_leaf_137_clk_regs sg13g2_dfrbpq_1
X_05586_ _02259_ VPWR _02261_ VGND _02257_ _02260_ sg13g2_o21ai_1
XFILLER_104_1014 VPWR VGND sg13g2_decap_8
X_07325_ _01461_ i_exotiny._1306_ _01598_ _02989_ VPWR VGND sg13g2_a21o_2
X_07256_ net2454 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[19\]
+ net1006 _00979_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_50_clk_regs clknet_5_14__leaf_clk_regs clknet_leaf_50_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06207_ net3188 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[15\]
+ net947 _00362_ VPWR VGND sg13g2_mux2_1
X_07187_ net1281 VPWR _02958_ VGND net3741 _02956_ sg13g2_o21ai_1
XFILLER_2_117 VPWR VGND sg13g2_fill_2
X_06138_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[29\]
+ net2389 net1046 _00307_ VPWR VGND sg13g2_mux2_1
XFILLER_105_557 VPWR VGND sg13g2_decap_8
X_08179__498 VPWR VGND net498 sg13g2_tiehi
X_06069_ VGND VPWR _01739_ _02516_ _00249_ _01388_ sg13g2_a21oi_1
XFILLER_87_964 VPWR VGND sg13g2_decap_8
XFILLER_101_763 VPWR VGND sg13g2_decap_4
XFILLER_100_262 VPWR VGND sg13g2_decap_8
XFILLER_73_124 VPWR VGND sg13g2_fill_1
XFILLER_46_338 VPWR VGND sg13g2_fill_2
XFILLER_27_530 VPWR VGND sg13g2_fill_2
XFILLER_42_511 VPWR VGND sg13g2_fill_2
XFILLER_11_953 VPWR VGND sg13g2_decap_8
X_08695__1293 VPWR VGND net1713 sg13g2_tiehi
X_09274__73 VPWR VGND net73 sg13g2_tiehi
XFILLER_7_968 VPWR VGND sg13g2_decap_8
XFILLER_9_1009 VPWR VGND sg13g2_decap_8
X_08590__1386 VPWR VGND net1806 sg13g2_tiehi
XFILLER_93_956 VPWR VGND sg13g2_decap_8
XFILLER_18_541 VPWR VGND sg13g2_fill_1
XFILLER_46_872 VPWR VGND sg13g2_fill_1
X_05440_ _02143_ _02144_ _02149_ VPWR VGND sg13g2_nor2_1
X_05371_ net1263 i_exotiny.i_wdg_top.do_cnt _02093_ VPWR VGND sg13g2_and2_1
X_09019__963 VPWR VGND net1383 sg13g2_tiehi
X_07110_ net1288 net1863 _00860_ VPWR VGND sg13g2_and2_1
X_08090_ net604 VGND VPWR _00171_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[27\]
+ clknet_leaf_85_clk_regs sg13g2_dfrbpq_1
Xclkload20 VPWR clkload20/Y clknet_leaf_32_clk_regs VGND sg13g2_inv_1
X_07041_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[11\]
+ net3109 net1013 _00802_ VPWR VGND sg13g2_mux2_1
Xclkload42 clknet_leaf_89_clk_regs clkload42/X VPWR VGND sg13g2_buf_8
Xclkload31 clkload31/Y clknet_leaf_145_clk_regs VPWR VGND sg13g2_inv_2
XFILLER_6_990 VPWR VGND sg13g2_decap_8
X_08992_ net1410 VGND VPWR net2011 i_exotiny._1160_\[13\] clknet_leaf_160_clk_regs
+ sg13g2_dfrbpq_1
X_08002__693 VPWR VGND net693 sg13g2_tiehi
X_09026__956 VPWR VGND net1376 sg13g2_tiehi
X_07943_ net87 VGND VPWR _00008_ i_exotiny._1737_ clknet_leaf_11_clk_regs sg13g2_dfrbpq_2
X_07874_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[12\]
+ net3473 net979 _01341_ VPWR VGND sg13g2_mux2_1
XFILLER_18_16 VPWR VGND sg13g2_fill_2
XFILLER_96_794 VPWR VGND sg13g2_fill_1
XFILLER_95_293 VPWR VGND sg13g2_decap_8
X_06825_ net3717 net1099 _02842_ VPWR VGND sg13g2_nor2_1
XFILLER_84_989 VPWR VGND sg13g2_decap_8
X_06756_ net1171 VPWR _02783_ VGND net3443 net1191 sg13g2_o21ai_1
XFILLER_70_149 VPWR VGND sg13g2_fill_1
X_06687_ _02724_ _02723_ net15 _02593_ net3551 VPWR VGND sg13g2_a22oi_1
X_05707_ net1918 net1058 _02351_ VPWR VGND sg13g2_nor2_1
XFILLER_51_330 VPWR VGND sg13g2_fill_1
X_09072__910 VPWR VGND net1330 sg13g2_tiehi
X_08962__1020 VPWR VGND net1440 sg13g2_tiehi
X_08426_ net259 VGND VPWR _00500_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[25\]
+ clknet_leaf_90_clk_regs sg13g2_dfrbpq_1
X_05638_ VGND VPWR net1061 _02299_ _00035_ _02297_ sg13g2_a21oi_1
Xclkload3 clknet_5_15__leaf_clk_regs clkload3/X VPWR VGND sg13g2_buf_8
X_08357_ net321 VGND VPWR net2674 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[27\]
+ clknet_leaf_98_clk_regs sg13g2_dfrbpq_1
X_09033__949 VPWR VGND net1369 sg13g2_tiehi
X_05569_ _01424_ VPWR _02249_ VGND i_exotiny._0315_\[7\] i_exotiny._0315_\[6\] sg13g2_o21ai_1
X_07308_ net2290 _02982_ net912 _01022_ VPWR VGND sg13g2_mux2_1
X_08288_ net390 VGND VPWR _00369_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[22\]
+ clknet_leaf_103_clk_regs sg13g2_dfrbpq_1
X_07239_ net3083 i_exotiny._0040_\[2\] net1004 _00962_ VPWR VGND sg13g2_mux2_1
XFILLER_106_811 VPWR VGND sg13g2_decap_8
XFILLER_105_354 VPWR VGND sg13g2_decap_8
XFILLER_106_888 VPWR VGND sg13g2_decap_8
Xfanout1205 net1206 net1205 VPWR VGND sg13g2_buf_8
Xfanout1227 _01378_ net1227 VPWR VGND sg13g2_buf_8
Xfanout1238 net1239 net1238 VPWR VGND sg13g2_buf_8
Xfanout1216 net1217 net1216 VPWR VGND sg13g2_buf_8
Xfanout1249 net3813 net1249 VPWR VGND sg13g2_buf_1
XFILLER_75_44 VPWR VGND sg13g2_fill_1
XFILLER_19_327 VPWR VGND sg13g2_fill_1
XFILLER_34_319 VPWR VGND sg13g2_fill_1
XFILLER_15_544 VPWR VGND sg13g2_fill_2
XFILLER_42_330 VPWR VGND sg13g2_fill_2
XFILLER_91_65 VPWR VGND sg13g2_fill_1
XFILLER_43_875 VPWR VGND sg13g2_fill_2
X_08782__1206 VPWR VGND net1626 sg13g2_tiehi
XFILLER_6_297 VPWR VGND sg13g2_fill_2
X_09049__934 VPWR VGND net1354 sg13g2_tiehi
XFILLER_66_912 VPWR VGND sg13g2_fill_1
XFILLER_27_4 VPWR VGND sg13g2_decap_8
X_04940_ _01644_ _01666_ _01629_ _01672_ VPWR VGND _01671_ sg13g2_nand4_1
XFILLER_93_720 VPWR VGND sg13g2_fill_1
X_04871_ _01381_ _01427_ net1248 _01603_ VPWR VGND sg13g2_nand3_1
X_07590_ net2028 _03163_ _03165_ VPWR VGND sg13g2_and2_1
X_06610_ i_exotiny._0314_\[16\] net1159 _02663_ VPWR VGND sg13g2_nor2_1
X_06541_ net2753 net881 _02620_ _02623_ VPWR VGND sg13g2_mux2_1
X_06472_ VGND VPWR net1166 _02615_ _02614_ net1139 sg13g2_a21oi_2
XFILLER_33_363 VPWR VGND sg13g2_fill_1
X_09260_ net241 VGND VPWR net2923 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[18\]
+ clknet_leaf_126_clk_regs sg13g2_dfrbpq_1
X_05423_ _01383_ _02131_ _02132_ VPWR VGND sg13g2_nor2_1
X_08211_ net466 VGND VPWR net2692 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[10\]
+ clknet_leaf_152_clk_regs sg13g2_dfrbpq_1
X_09191_ net790 VGND VPWR net2242 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[13\]
+ clknet_leaf_78_clk_regs sg13g2_dfrbpq_1
X_08758__1230 VPWR VGND net1650 sg13g2_tiehi
X_05354_ _02076_ net3326 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set[0]
+ VPWR VGND sg13g2_nand2b_1
X_08142_ net543 VGND VPWR _00223_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[6\]
+ clknet_leaf_155_clk_regs sg13g2_dfrbpq_1
X_08073_ net621 VGND VPWR net2970 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[10\]
+ clknet_leaf_85_clk_regs sg13g2_dfrbpq_1
Xclkbuf_5_24__f_clk_regs clknet_4_12_0_clk_regs clknet_5_24__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_05285_ _02010_ VPWR _02011_ VGND i_exotiny._0036_\[0\] _01755_ sg13g2_o21ai_1
XFILLER_106_118 VPWR VGND sg13g2_decap_8
X_07024_ net3320 net887 _02928_ _02930_ VPWR VGND sg13g2_mux2_1
XFILLER_1_908 VPWR VGND sg13g2_decap_8
XFILLER_103_825 VPWR VGND sg13g2_decap_8
XFILLER_88_547 VPWR VGND sg13g2_fill_1
X_08975_ net1427 VGND VPWR net3740 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[0\]
+ clknet_leaf_165_clk_regs sg13g2_dfrbpq_2
Xhold37 i_exotiny.i_wb_spi.state_r\[30\] VPWR VGND net1864 sg13g2_dlygate4sd3_1
XFILLER_102_357 VPWR VGND sg13g2_decap_8
Xhold26 i_exotiny.i_wb_spi.state_r\[10\] VPWR VGND net1853 sg13g2_dlygate4sd3_1
Xhold15 _00874_ VPWR VGND net1842 sg13g2_dlygate4sd3_1
X_07926_ net722 VGND VPWR net1948 i_exotiny._1924_\[19\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
XFILLER_60_1001 VPWR VGND sg13g2_fill_1
Xhold1911 i_exotiny._1611_\[14\] VPWR VGND net3738 sg13g2_dlygate4sd3_1
Xhold1900 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[2\]
+ VPWR VGND net3727 sg13g2_dlygate4sd3_1
Xhold59 _03157_ VPWR VGND net1886 sg13g2_dlygate4sd3_1
Xhold48 i_exotiny.i_wdg_top.o_wb_dat\[12\] VPWR VGND net1875 sg13g2_dlygate4sd3_1
XFILLER_56_422 VPWR VGND sg13g2_fill_1
XFILLER_28_102 VPWR VGND sg13g2_fill_2
Xhold1922 i_exotiny._0369_\[13\] VPWR VGND net3749 sg13g2_dlygate4sd3_1
Xhold1933 _00513_ VPWR VGND net3760 sg13g2_dlygate4sd3_1
Xhold1944 _03011_ VPWR VGND net3771 sg13g2_dlygate4sd3_1
Xhold1955 i_exotiny._2055_\[0\] VPWR VGND net3782 sg13g2_dlygate4sd3_1
Xhold1966 _00075_ VPWR VGND net3793 sg13g2_dlygate4sd3_1
XFILLER_56_444 VPWR VGND sg13g2_decap_8
Xhold1988 i_exotiny._1660_ VPWR VGND net3815 sg13g2_dlygate4sd3_1
X_07857_ _03226_ net2121 net984 _01327_ VPWR VGND sg13g2_mux2_1
Xhold1977 i_exotiny._0077_\[0\] VPWR VGND net3804 sg13g2_dlygate4sd3_1
XFILLER_71_414 VPWR VGND sg13g2_fill_2
X_06808_ VGND VPWR net1096 net3698 _00677_ _02827_ sg13g2_a21oi_1
X_07788_ net3525 net3481 net892 _01267_ VPWR VGND sg13g2_mux2_1
Xhold1999 i_exotiny._0079_\[2\] VPWR VGND net3826 sg13g2_dlygate4sd3_1
X_06739_ _02768_ VPWR _02769_ VGND i_exotiny._0369_\[7\] net1192 sg13g2_o21ai_1
X_08903__1079 VPWR VGND net1499 sg13g2_tiehi
XFILLER_52_650 VPWR VGND sg13g2_decap_8
XFILLER_25_864 VPWR VGND sg13g2_fill_1
XFILLER_24_396 VPWR VGND sg13g2_fill_2
X_08409_ net276 VGND VPWR net2930 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[8\]
+ clknet_leaf_93_clk_regs sg13g2_dfrbpq_1
XFILLER_4_724 VPWR VGND sg13g2_fill_1
X_08124__570 VPWR VGND net570 sg13g2_tiehi
XFILLER_106_685 VPWR VGND sg13g2_decap_8
XFILLER_105_151 VPWR VGND sg13g2_decap_8
Xfanout1013 net1014 net1013 VPWR VGND sg13g2_buf_8
Xfanout1002 _03194_ net1002 VPWR VGND sg13g2_buf_8
Xfanout1024 _02615_ net1024 VPWR VGND sg13g2_buf_8
XFILLER_67_709 VPWR VGND sg13g2_fill_1
XFILLER_0_952 VPWR VGND sg13g2_decap_8
Xfanout1035 net1036 net1035 VPWR VGND sg13g2_buf_8
Xfanout1046 net1047 net1046 VPWR VGND sg13g2_buf_8
X_09009__973 VPWR VGND net1393 sg13g2_tiehi
Xfanout1057 _02424_ net1057 VPWR VGND sg13g2_buf_8
X_08548__108 VPWR VGND net108 sg13g2_tiehi
Xfanout1068 _02718_ net1068 VPWR VGND sg13g2_buf_8
Xfanout1079 net1085 net1079 VPWR VGND sg13g2_buf_8
X_08836__1152 VPWR VGND net1572 sg13g2_tiehi
XFILLER_35_606 VPWR VGND sg13g2_fill_1
XFILLER_47_499 VPWR VGND sg13g2_fill_1
XFILLER_74_285 VPWR VGND sg13g2_fill_2
XFILLER_34_138 VPWR VGND sg13g2_fill_2
X_09016__966 VPWR VGND net1386 sg13g2_tiehi
Xclkbuf_leaf_178_clk_regs clknet_5_1__leaf_clk_regs clknet_leaf_178_clk_regs VPWR
+ VGND sg13g2_buf_8
Xclkbuf_leaf_107_clk_regs clknet_5_28__leaf_clk_regs clknet_leaf_107_clk_regs VPWR
+ VGND sg13g2_buf_8
Xhold518 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[23\]
+ VPWR VGND net2345 sg13g2_dlygate4sd3_1
Xhold507 _00305_ VPWR VGND net2334 sg13g2_dlygate4sd3_1
Xhold529 _00755_ VPWR VGND net2356 sg13g2_dlygate4sd3_1
X_05070_ _01799_ _01801_ _01802_ VPWR VGND sg13g2_nor2_1
XFILLER_98_867 VPWR VGND sg13g2_decap_8
X_09062__920 VPWR VGND net1340 sg13g2_tiehi
XFILLER_97_366 VPWR VGND sg13g2_decap_8
Xhold1207 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[14\]
+ VPWR VGND net3034 sg13g2_dlygate4sd3_1
X_08760_ net1648 VGND VPWR net2556 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[23\]
+ clknet_leaf_87_clk_regs sg13g2_dfrbpq_1
Xhold1218 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[18\]
+ VPWR VGND net3045 sg13g2_dlygate4sd3_1
X_05972_ _02420_ _02492_ _02493_ VPWR VGND sg13g2_nor2_2
Xhold1229 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[26\]
+ VPWR VGND net3056 sg13g2_dlygate4sd3_1
X_08691_ net1717 VGND VPWR _00749_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[18\]
+ clknet_leaf_103_clk_regs sg13g2_dfrbpq_1
X_04923_ net1223 _01613_ _01623_ _01655_ VPWR VGND sg13g2_nor3_2
X_09023__959 VPWR VGND net1379 sg13g2_tiehi
X_07711_ net2335 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[8\]
+ net993 _01207_ VPWR VGND sg13g2_mux2_1
XFILLER_18_0 VPWR VGND sg13g2_fill_2
X_04854_ _01590_ i_exotiny.i_wb_spi.cnt_presc_r\[4\] _01573_ VPWR VGND sg13g2_xnor2_1
X_07642_ net2706 net2952 net896 _01150_ VPWR VGND sg13g2_mux2_1
Xclkbuf_5_8__f_clk_regs clknet_4_4_0_clk_regs clknet_5_8__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07573_ net3201 net1830 _03154_ VPWR VGND sg13g2_and2_1
X_04785_ _01535_ net1230 _01534_ VPWR VGND sg13g2_xnor2_1
X_06524_ net3132 net3054 net932 _00599_ VPWR VGND sg13g2_mux2_1
XFILLER_33_160 VPWR VGND sg13g2_fill_1
X_06455_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[24\]
+ net3068 net938 _00542_ VPWR VGND sg13g2_mux2_1
X_09243_ net564 VGND VPWR net3492 i_exotiny._0022_\[1\] clknet_leaf_127_clk_regs sg13g2_dfrbpq_2
X_05406_ _02119_ i_exotiny._2034_\[5\] i_exotiny._2034_\[6\] _02115_ VPWR VGND sg13g2_and3_1
X_09174_ net808 VGND VPWR _01229_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[30\]
+ clknet_leaf_172_clk_regs sg13g2_dfrbpq_1
XFILLER_21_366 VPWR VGND sg13g2_fill_1
X_06386_ VGND VPWR net3647 _02180_ _02575_ _02574_ sg13g2_a21oi_1
X_08125_ net569 VGND VPWR _00206_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[30\]
+ clknet_leaf_121_clk_regs sg13g2_dfrbpq_1
X_05337_ _01912_ VPWR _02061_ VGND _02059_ _02060_ sg13g2_o21ai_1
X_08056_ net638 VGND VPWR _00137_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[25\]
+ clknet_leaf_55_clk_regs sg13g2_dfrbpq_1
X_05268_ _01994_ _01786_ i_exotiny._0017_\[0\] _01769_ i_exotiny._0022_\[0\] VPWR
+ VGND sg13g2_a22oi_1
Xoutput38 net38 uo_out[4] VPWR VGND sg13g2_buf_1
Xoutput27 net27 uio_out[1] VPWR VGND sg13g2_buf_1
X_07007_ net2972 net3130 net918 _00774_ VPWR VGND sg13g2_mux2_1
X_05199_ _01927_ _01779_ i_exotiny._0020_\[1\] _01773_ i_exotiny._0019_\[1\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_103_677 VPWR VGND sg13g2_fill_1
XFILLER_103_666 VPWR VGND sg13g2_decap_8
X_08958_ net1444 VGND VPWR net2663 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[24\]
+ clknet_leaf_75_clk_regs sg13g2_dfrbpq_1
XFILLER_76_528 VPWR VGND sg13g2_fill_1
XFILLER_5_1001 VPWR VGND sg13g2_decap_8
Xhold1752 _03171_ VPWR VGND net3579 sg13g2_dlygate4sd3_1
Xhold1741 _00024_ VPWR VGND net3568 sg13g2_dlygate4sd3_1
X_08889_ net1513 VGND VPWR _00947_ i_exotiny.i_wb_spi.dat_rx_r\[19\] clknet_leaf_63_clk_regs
+ sg13g2_dfrbpq_1
X_07909_ net739 VGND VPWR net1979 i_exotiny._1924_\[2\] clknet_leaf_31_clk_regs sg13g2_dfrbpq_1
Xhold1730 _00932_ VPWR VGND net3557 sg13g2_dlygate4sd3_1
XFILLER_71_200 VPWR VGND sg13g2_fill_1
Xhold1763 _00929_ VPWR VGND net3590 sg13g2_dlygate4sd3_1
Xhold1796 i_exotiny.i_wb_spi.dat_rx_r\[28\] VPWR VGND net3623 sg13g2_dlygate4sd3_1
Xhold1774 i_exotiny._0369_\[29\] VPWR VGND net3601 sg13g2_dlygate4sd3_1
Xhold1785 i_exotiny._0315_\[15\] VPWR VGND net3612 sg13g2_dlygate4sd3_1
XFILLER_71_233 VPWR VGND sg13g2_fill_1
XFILLER_16_127 VPWR VGND sg13g2_fill_1
XFILLER_44_458 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_5_clk_regs clknet_5_3__leaf_clk_regs clknet_leaf_5_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08478__202 VPWR VGND net202 sg13g2_tiehi
XFILLER_4_532 VPWR VGND sg13g2_fill_1
XFILLER_106_482 VPWR VGND sg13g2_decap_8
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_06240_ net3334 net3087 net1038 _00389_ VPWR VGND sg13g2_mux2_1
X_06171_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[19\]
+ net2238 net950 _00333_ VPWR VGND sg13g2_mux2_1
XFILLER_105_909 VPWR VGND sg13g2_decap_8
Xhold326 _00092_ VPWR VGND net2153 sg13g2_dlygate4sd3_1
Xhold304 _01153_ VPWR VGND net2131 sg13g2_dlygate4sd3_1
X_05122_ _01852_ _01772_ i_exotiny._0033_\[2\] _01760_ i_exotiny._0014_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold315 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[14\]
+ VPWR VGND net2142 sg13g2_dlygate4sd3_1
Xhold337 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[25\]
+ VPWR VGND net2164 sg13g2_dlygate4sd3_1
Xhold348 _00891_ VPWR VGND net2175 sg13g2_dlygate4sd3_1
Xhold359 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[5\]
+ VPWR VGND net2186 sg13g2_dlygate4sd3_1
X_05053_ net1236 _01759_ _01762_ _01785_ VPWR VGND sg13g2_nor3_2
X_08138__547 VPWR VGND net547 sg13g2_tiehi
Xhold1004 _00815_ VPWR VGND net2831 sg13g2_dlygate4sd3_1
X_08812_ net1596 VGND VPWR _00870_ i_exotiny.i_wb_spi.state_r\[11\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_75_clk_regs clknet_5_26__leaf_clk_regs clknet_leaf_75_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold1015 _01090_ VPWR VGND net2842 sg13g2_dlygate4sd3_1
Xhold1026 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[31\]
+ VPWR VGND net2853 sg13g2_dlygate4sd3_1
X_05955_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[20\]
+ net2234 net968 _00164_ VPWR VGND sg13g2_mux2_1
X_08743_ net1665 VGND VPWR net2921 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[6\]
+ clknet_leaf_84_clk_regs sg13g2_dfrbpq_1
Xhold1048 _00598_ VPWR VGND net2875 sg13g2_dlygate4sd3_1
Xhold1037 i_exotiny._0314_\[17\] VPWR VGND net2864 sg13g2_dlygate4sd3_1
Xhold1059 i_exotiny._0314_\[30\] VPWR VGND net2886 sg13g2_dlygate4sd3_1
XFILLER_38_241 VPWR VGND sg13g2_fill_1
XFILLER_39_786 VPWR VGND sg13g2_fill_2
X_04906_ net1222 _01616_ _01620_ _01638_ VPWR VGND sg13g2_nor3_2
XFILLER_94_892 VPWR VGND sg13g2_decap_8
XFILLER_54_734 VPWR VGND sg13g2_fill_1
X_08674_ net1734 VGND VPWR net2678 i_exotiny._0034_\[1\] clknet_leaf_111_clk_regs
+ sg13g2_dfrbpq_2
X_08114__580 VPWR VGND net580 sg13g2_tiehi
X_05886_ _01470_ _02465_ _02470_ _02472_ VPWR VGND sg13g2_nor3_2
XFILLER_38_285 VPWR VGND sg13g2_fill_2
X_04837_ _01571_ _01576_ _01577_ VPWR VGND sg13g2_nor2b_2
X_07625_ _02477_ _02517_ _03187_ VPWR VGND sg13g2_nor2_2
XFILLER_42_929 VPWR VGND sg13g2_fill_2
X_07556_ _03134_ VPWR _03143_ VGND net3681 _03140_ sg13g2_o21ai_1
X_04768_ net1193 net1169 _01518_ _01519_ VPWR VGND sg13g2_nor3_2
X_06507_ i_exotiny._0041_\[3\] net874 _02614_ _02619_ VPWR VGND sg13g2_mux2_1
X_09226_ net753 VGND VPWR net2870 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[16\]
+ clknet_leaf_136_clk_regs sg13g2_dfrbpq_1
X_04699_ net1251 _01456_ _01457_ VPWR VGND sg13g2_nor2_1
X_07487_ VGND VPWR _01390_ net903 _01073_ _03110_ sg13g2_a21oi_1
XFILLER_21_196 VPWR VGND sg13g2_fill_2
X_06438_ net3344 i_exotiny._0039_\[3\] net934 _00525_ VPWR VGND sg13g2_mux2_1
X_06369_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[28\]
+ net2995 net1028 _00499_ VPWR VGND sg13g2_mux2_1
X_09157_ net825 VGND VPWR net2580 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[13\]
+ clknet_leaf_173_clk_regs sg13g2_dfrbpq_1
X_08108_ net586 VGND VPWR net2596 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[13\]
+ clknet_leaf_125_clk_regs sg13g2_dfrbpq_1
X_09088_ net1314 VGND VPWR _01143_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[8\]
+ clknet_leaf_141_clk_regs sg13g2_dfrbpq_1
X_08039_ net655 VGND VPWR net2932 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[8\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
X_08121__573 VPWR VGND net573 sg13g2_tiehi
Xhold871 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[20\]
+ VPWR VGND net2698 sg13g2_dlygate4sd3_1
Xhold860 _01145_ VPWR VGND net2687 sg13g2_dlygate4sd3_1
Xhold882 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[24\]
+ VPWR VGND net2709 sg13g2_dlygate4sd3_1
XFILLER_103_430 VPWR VGND sg13g2_decap_8
Xhold893 i_exotiny._0029_\[3\] VPWR VGND net2720 sg13g2_dlygate4sd3_1
XFILLER_104_986 VPWR VGND sg13g2_decap_8
Xhold1571 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[26\]
+ VPWR VGND net3398 sg13g2_dlygate4sd3_1
X_09006__976 VPWR VGND net1396 sg13g2_tiehi
Xhold1560 i_exotiny._1840_\[11\] VPWR VGND net3387 sg13g2_dlygate4sd3_1
Xhold1582 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[25\]
+ VPWR VGND net3409 sg13g2_dlygate4sd3_1
XFILLER_84_380 VPWR VGND sg13g2_fill_2
Xhold1593 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[23\]
+ VPWR VGND net3420 sg13g2_dlygate4sd3_1
XFILLER_44_255 VPWR VGND sg13g2_fill_1
XFILLER_16_93 VPWR VGND sg13g2_fill_1
X_09052__930 VPWR VGND net1350 sg13g2_tiehi
X_08640__1337 VPWR VGND net1757 sg13g2_tiehi
X_09013__969 VPWR VGND net1389 sg13g2_tiehi
XFILLER_5_896 VPWR VGND sg13g2_decap_8
XFILLER_80_1026 VPWR VGND sg13g2_fill_2
X_08567__70 VPWR VGND net70 sg13g2_tiehi
XFILLER_83_807 VPWR VGND sg13g2_fill_2
X_05740_ _02368_ net3703 _02377_ VPWR VGND sg13g2_xor2_1
X_05671_ net1947 net1062 _02324_ VPWR VGND sg13g2_nor2_1
XFILLER_24_929 VPWR VGND sg13g2_fill_1
X_04622_ _01384_ net1232 VPWR VGND sg13g2_inv_2
X_08390_ net288 VGND VPWR _00471_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[28\]
+ clknet_leaf_139_clk_regs sg13g2_dfrbpq_1
X_07410_ net1080 _03058_ _03059_ _03060_ VPWR VGND sg13g2_nor3_1
X_07341_ _02993_ _02996_ _03003_ _03005_ VPWR VGND sg13g2_nor3_1
Xclkbuf_leaf_122_clk_regs clknet_5_22__leaf_clk_regs clknet_leaf_122_clk_regs VPWR
+ VGND sg13g2_buf_8
X_07272_ _02977_ net3173 net1006 _00991_ VPWR VGND sg13g2_mux2_1
X_06223_ _02543_ net2305 net945 _00376_ VPWR VGND sg13g2_mux2_1
X_09168__814 VPWR VGND net814 sg13g2_tiehi
X_09011_ net1391 VGND VPWR net3581 i_exotiny._0079_\[4\] clknet_leaf_160_clk_regs
+ sg13g2_dfrbpq_1
X_06154_ i_exotiny._0028_\[2\] net2166 net952 _00316_ VPWR VGND sg13g2_mux2_1
Xhold101 i_exotiny.i_wb_spi.spi_sdo_o VPWR VGND net1928 sg13g2_dlygate4sd3_1
XFILLER_105_706 VPWR VGND sg13g2_decap_8
Xhold112 i_exotiny._1924_\[14\] VPWR VGND net1939 sg13g2_dlygate4sd3_1
Xhold134 i_exotiny._1924_\[1\] VPWR VGND net1961 sg13g2_dlygate4sd3_1
X_05105_ _01832_ _01833_ _01828_ _01835_ VPWR VGND sg13g2_nand3_1
Xhold123 _01040_ VPWR VGND net1950 sg13g2_dlygate4sd3_1
XFILLER_99_940 VPWR VGND sg13g2_decap_8
Xhold145 i_exotiny.i_wb_spi.cnt_hbit_r\[4\] VPWR VGND net1972 sg13g2_dlygate4sd3_1
X_06085_ net2761 net3366 net960 _00261_ VPWR VGND sg13g2_mux2_1
Xhold156 _00051_ VPWR VGND net1983 sg13g2_dlygate4sd3_1
Xhold167 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[21\]
+ VPWR VGND net1994 sg13g2_dlygate4sd3_1
Xhold178 _00041_ VPWR VGND net2005 sg13g2_dlygate4sd3_1
Xhold189 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[26\]
+ VPWR VGND net2016 sg13g2_dlygate4sd3_1
X_05036_ i_exotiny._0079_\[2\] i_exotiny._0079_\[3\] net1221 _01768_ VPWR VGND sg13g2_or3_1
XFILLER_101_934 VPWR VGND sg13g2_decap_8
XFILLER_100_444 VPWR VGND sg13g2_decap_8
XFILLER_85_155 VPWR VGND sg13g2_fill_1
X_08468__212 VPWR VGND net212 sg13g2_tiehi
X_06987_ net2355 _02924_ net1021 _00759_ VPWR VGND sg13g2_mux2_1
X_05938_ i_exotiny._0020_\[3\] net3081 net966 _00147_ VPWR VGND sg13g2_mux2_1
X_09175__807 VPWR VGND net807 sg13g2_tiehi
XFILLER_37_59 VPWR VGND sg13g2_fill_1
X_08726_ net1682 VGND VPWR _00784_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[21\]
+ clknet_leaf_120_clk_regs sg13g2_dfrbpq_1
X_08657_ net1740 VGND VPWR net2928 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[26\]
+ clknet_leaf_149_clk_regs sg13g2_dfrbpq_1
X_05869_ VGND VPWR _01911_ _02267_ _02456_ _02428_ sg13g2_a21oi_1
X_07608_ net3722 _03175_ _03176_ VPWR VGND sg13g2_and2_1
X_08588_ net1808 VGND VPWR net3633 i_exotiny._6090_\[0\] clknet_leaf_9_clk_regs sg13g2_dfrbpq_1
X_07539_ _03126_ _03131_ _01443_ _03132_ VPWR VGND sg13g2_nand3_1
X_09209_ net770 VGND VPWR net2854 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[31\]
+ clknet_leaf_76_clk_regs sg13g2_dfrbpq_1
X_08475__205 VPWR VGND net205 sg13g2_tiehi
XFILLER_10_689 VPWR VGND sg13g2_fill_2
Xhold690 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[30\]
+ VPWR VGND net2517 sg13g2_dlygate4sd3_1
XFILLER_1_343 VPWR VGND sg13g2_fill_2
XFILLER_2_866 VPWR VGND sg13g2_decap_8
XFILLER_104_783 VPWR VGND sg13g2_decap_8
X_08195__482 VPWR VGND net482 sg13g2_tiehi
XFILLER_76_100 VPWR VGND sg13g2_fill_1
X_08658__1319 VPWR VGND net1739 sg13g2_tiehi
XFILLER_76_177 VPWR VGND sg13g2_fill_2
XFILLER_18_734 VPWR VGND sg13g2_fill_1
Xhold1390 _00741_ VPWR VGND net3217 sg13g2_dlygate4sd3_1
XFILLER_17_255 VPWR VGND sg13g2_fill_2
XFILLER_27_70 VPWR VGND sg13g2_fill_2
XFILLER_45_553 VPWR VGND sg13g2_fill_1
XFILLER_14_995 VPWR VGND sg13g2_fill_2
XFILLER_40_280 VPWR VGND sg13g2_fill_2
XFILLER_43_91 VPWR VGND sg13g2_fill_2
X_08916__1066 VPWR VGND net1486 sg13g2_tiehi
X_10679_ _10679_/A net32 VPWR VGND sg13g2_buf_1
X_08104__590 VPWR VGND net590 sg13g2_tiehi
XFILLER_99_269 VPWR VGND sg13g2_decap_8
XFILLER_101_219 VPWR VGND sg13g2_decap_8
XFILLER_96_921 VPWR VGND sg13g2_decap_8
X_06910_ i_exotiny.i_rstctl.cnt\[1\] i_exotiny.i_rstctl.cnt\[5\] net1883 _02910_ VPWR
+ VGND i_exotiny.i_rstctl.cnt\[4\] sg13g2_nand4_1
XFILLER_67_100 VPWR VGND sg13g2_fill_1
X_07890_ net2534 net886 _03228_ _03230_ VPWR VGND sg13g2_mux2_1
XFILLER_96_998 VPWR VGND sg13g2_decap_8
X_06841_ net1128 _02853_ _02854_ _02855_ VPWR VGND sg13g2_nor3_1
XFILLER_83_626 VPWR VGND sg13g2_fill_1
X_06772_ VGND VPWR _02794_ _02796_ _02797_ net1135 sg13g2_a21oi_1
XFILLER_55_328 VPWR VGND sg13g2_fill_1
X_08511_ net169 VGND VPWR net3118 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[31\]
+ clknet_leaf_109_clk_regs sg13g2_dfrbpq_1
X_05723_ net1114 i_exotiny._1924_\[31\] _02363_ VPWR VGND sg13g2_nor2b_1
X_08627__742 VPWR VGND net742 sg13g2_tiehi
X_08442_ net242 VGND VPWR _00516_ i_exotiny._2025_\[4\] clknet_leaf_29_clk_regs sg13g2_dfrbpq_2
X_05654_ VGND VPWR net1067 _02311_ _00039_ _02309_ sg13g2_a21oi_1
X_08111__583 VPWR VGND net583 sg13g2_tiehi
X_04605_ VPWR _01367_ i_exotiny._1615_\[1\] VGND sg13g2_inv_1
X_08373_ net305 VGND VPWR net2827 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[11\]
+ clknet_leaf_133_clk_regs sg13g2_dfrbpq_1
X_05585_ _02260_ i_exotiny._1306_ i_exotiny._0352_ VPWR VGND sg13g2_nand2_1
X_07324_ VGND VPWR i_exotiny._1306_ _01461_ _02988_ _01598_ sg13g2_a21oi_1
X_07255_ net2616 net2339 net1003 _00978_ VPWR VGND sg13g2_mux2_1
X_06206_ net2566 net2794 net948 _00361_ VPWR VGND sg13g2_mux2_1
X_07186_ VGND VPWR _01361_ _02956_ _00925_ net3773 sg13g2_a21oi_1
XFILLER_105_536 VPWR VGND sg13g2_decap_8
X_09181__800 VPWR VGND net800 sg13g2_tiehi
Xclkbuf_leaf_90_clk_regs clknet_5_31__leaf_clk_regs clknet_leaf_90_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06137_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[28\]
+ net2709 net1043 _00306_ VPWR VGND sg13g2_mux2_1
X_06068_ _02516_ net2140 _01701_ VPWR VGND sg13g2_nand2_1
X_05019_ VGND VPWR net1267 i_exotiny._6090_\[3\] _01751_ _01750_ sg13g2_a21oi_1
XFILLER_86_431 VPWR VGND sg13g2_fill_1
XFILLER_100_241 VPWR VGND sg13g2_decap_8
X_09042__940 VPWR VGND net1360 sg13g2_tiehi
XFILLER_39_380 VPWR VGND sg13g2_fill_1
XFILLER_104_75 VPWR VGND sg13g2_fill_1
XFILLER_104_64 VPWR VGND sg13g2_fill_1
X_09003__979 VPWR VGND net1399 sg13g2_tiehi
X_08709_ net1699 VGND VPWR _00767_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[4\]
+ clknet_leaf_120_clk_regs sg13g2_dfrbpq_1
XFILLER_42_578 VPWR VGND sg13g2_decap_4
XFILLER_42_589 VPWR VGND sg13g2_fill_2
XFILLER_6_402 VPWR VGND sg13g2_fill_1
XFILLER_7_947 VPWR VGND sg13g2_decap_8
XFILLER_6_435 VPWR VGND sg13g2_fill_1
X_09227__752 VPWR VGND net752 sg13g2_tiehi
XFILLER_104_580 VPWR VGND sg13g2_fill_2
X_08607__1369 VPWR VGND net1789 sg13g2_tiehi
XFILLER_93_935 VPWR VGND sg13g2_decap_8
XFILLER_77_497 VPWR VGND sg13g2_fill_2
XFILLER_38_80 VPWR VGND sg13g2_decap_8
XFILLER_80_607 VPWR VGND sg13g2_fill_1
X_09158__824 VPWR VGND net824 sg13g2_tiehi
XFILLER_45_350 VPWR VGND sg13g2_fill_2
X_09234__745 VPWR VGND net745 sg13g2_tiehi
XFILLER_33_578 VPWR VGND sg13g2_fill_2
X_05370_ net1832 _02076_ net1112 _02092_ VPWR VGND sg13g2_nor3_1
XFILLER_14_792 VPWR VGND sg13g2_fill_2
XFILLER_9_240 VPWR VGND sg13g2_fill_2
X_08458__222 VPWR VGND net222 sg13g2_tiehi
Xclkload10 clknet_leaf_6_clk_regs clkload10/Y VPWR VGND sg13g2_inv_4
Xclkbuf_5_23__f_clk_regs clknet_4_11_0_clk_regs clknet_5_23__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07040_ net2920 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[6\]
+ net1017 _00801_ VPWR VGND sg13g2_mux2_1
Xclkload43 VPWR clkload43/Y clknet_leaf_91_clk_regs VGND sg13g2_inv_1
Xclkload21 clknet_leaf_26_clk_regs clkload21/Y VPWR VGND sg13g2_inv_4
Xclkload32 clknet_leaf_138_clk_regs clkload32/Y VPWR VGND sg13g2_inv_4
X_09165__817 VPWR VGND net817 sg13g2_tiehi
XFILLER_48_0 VPWR VGND sg13g2_fill_2
XFILLER_88_718 VPWR VGND sg13g2_fill_2
X_08991_ net1411 VGND VPWR net2078 i_exotiny._1160_\[12\] clknet_leaf_18_clk_regs
+ sg13g2_dfrbpq_1
X_07942_ net86 VGND VPWR net3522 i_exotiny._1715_ clknet_leaf_27_clk_regs sg13g2_dfrbpq_2
X_07873_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[11\]
+ net2188 net980 _01340_ VPWR VGND sg13g2_mux2_1
XFILLER_95_272 VPWR VGND sg13g2_decap_8
XFILLER_84_946 VPWR VGND sg13g2_fill_2
X_06824_ VGND VPWR net3501 net1134 _02841_ _02840_ sg13g2_a21oi_1
X_08465__215 VPWR VGND net215 sg13g2_tiehi
X_06755_ _02782_ VPWR _00669_ VGND net1137 _02781_ sg13g2_o21ai_1
X_05706_ VGND VPWR net1058 _02349_ _00052_ _02350_ sg13g2_a21oi_1
X_06686_ _02723_ _01390_ net1233 _01391_ VPWR VGND sg13g2_and3_2
XFILLER_24_545 VPWR VGND sg13g2_fill_1
XFILLER_36_383 VPWR VGND sg13g2_fill_2
X_08425_ net260 VGND VPWR net2996 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[24\]
+ clknet_leaf_91_clk_regs sg13g2_dfrbpq_1
X_05637_ VGND VPWR i_exotiny._1615_\[1\] net1119 _02299_ _02298_ sg13g2_a21oi_1
X_08356_ net322 VGND VPWR net3207 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[26\]
+ clknet_leaf_107_clk_regs sg13g2_dfrbpq_1
X_08185__492 VPWR VGND net492 sg13g2_tiehi
X_07307_ net880 net3168 _02978_ _02982_ VPWR VGND sg13g2_mux2_1
Xclkload4 clknet_5_23__leaf_clk_regs clkload4/X VPWR VGND sg13g2_buf_8
X_05568_ VGND VPWR _01385_ _02246_ i_exotiny._1489_\[1\] net3678 sg13g2_a21oi_1
X_08287_ net391 VGND VPWR net2370 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[21\]
+ clknet_leaf_107_clk_regs sg13g2_dfrbpq_1
X_05499_ _02194_ net3737 net1069 VPWR VGND sg13g2_nand2_1
X_07238_ net2889 i_exotiny._0040_\[1\] net1005 _00961_ VPWR VGND sg13g2_mux2_1
X_08472__208 VPWR VGND net208 sg13g2_tiehi
X_07169_ net2861 net2608 net1010 _00917_ VPWR VGND sg13g2_mux2_1
XFILLER_4_939 VPWR VGND sg13g2_decap_8
XFILLER_106_867 VPWR VGND sg13g2_decap_8
XFILLER_105_333 VPWR VGND sg13g2_decap_8
Xfanout1228 net3839 net1228 VPWR VGND sg13g2_buf_8
Xfanout1206 _02256_ net1206 VPWR VGND sg13g2_buf_2
XFILLER_8_1021 VPWR VGND sg13g2_decap_8
Xfanout1217 _01503_ net1217 VPWR VGND sg13g2_buf_8
X_08192__485 VPWR VGND net485 sg13g2_tiehi
Xfanout1239 net3836 net1239 VPWR VGND sg13g2_buf_2
XFILLER_28_862 VPWR VGND sg13g2_fill_1
XFILLER_43_887 VPWR VGND sg13g2_fill_2
XFILLER_7_733 VPWR VGND sg13g2_fill_2
X_08101__593 VPWR VGND net593 sg13g2_tiehi
XFILLER_65_423 VPWR VGND sg13g2_decap_8
X_09258__509 VPWR VGND net509 sg13g2_tiehi
XFILLER_1_42 VPWR VGND sg13g2_decap_8
X_04870_ net1271 net1266 net1268 _01602_ VPWR VGND sg13g2_or3_1
XFILLER_37_147 VPWR VGND sg13g2_fill_1
Xclkbuf_5_7__f_clk_regs clknet_4_3_0_clk_regs clknet_5_7__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_53_607 VPWR VGND sg13g2_fill_2
X_06540_ net2617 _02622_ net932 _00614_ VPWR VGND sg13g2_mux2_1
X_06471_ _02419_ _02518_ _02614_ VPWR VGND sg13g2_nor2_2
X_05422_ _01536_ _02130_ net1146 _02131_ VPWR VGND sg13g2_nand3_1
X_08210_ net467 VGND VPWR _00291_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[9\]
+ clknet_leaf_153_clk_regs sg13g2_dfrbpq_1
X_09190_ net791 VGND VPWR _01245_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[12\]
+ clknet_leaf_77_clk_regs sg13g2_dfrbpq_1
XFILLER_60_194 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_29_clk_regs clknet_5_8__leaf_clk_regs clknet_leaf_29_clk_regs VPWR VGND
+ sg13g2_buf_8
X_05353_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set[0]
+ _02074_ _02075_ VPWR VGND sg13g2_nor2_1
XFILLER_14_1026 VPWR VGND sg13g2_fill_2
X_08141_ net544 VGND VPWR _00222_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[5\]
+ clknet_leaf_132_clk_regs sg13g2_dfrbpq_1
XFILLER_101_1018 VPWR VGND sg13g2_decap_8
X_08072_ net622 VGND VPWR _00153_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[9\]
+ clknet_leaf_92_clk_regs sg13g2_dfrbpq_1
X_09032__950 VPWR VGND net1370 sg13g2_tiehi
X_05284_ _02004_ _02009_ _02000_ _02010_ VPWR VGND sg13g2_nand3_1
X_07023_ net3183 net3301 net918 _00790_ VPWR VGND sg13g2_mux2_1
X_08653__1324 VPWR VGND net1744 sg13g2_tiehi
XFILLER_103_804 VPWR VGND sg13g2_decap_8
XFILLER_88_504 VPWR VGND sg13g2_fill_2
XFILLER_102_336 VPWR VGND sg13g2_decap_8
X_08974_ net1428 VGND VPWR _01032_ i_exotiny._0550_ clknet_leaf_14_clk_regs sg13g2_dfrbpq_2
Xhold27 i_exotiny.i_wb_spi.state_r\[31\] VPWR VGND net1854 sg13g2_dlygate4sd3_1
Xhold38 i_exotiny.i_wb_spi.state_r\[18\] VPWR VGND net1865 sg13g2_dlygate4sd3_1
Xhold16 i_exotiny.i_wb_spi.state_r\[25\] VPWR VGND net1843 sg13g2_dlygate4sd3_1
Xhold1901 i_exotiny.i_wb_spi.cnt_presc_r\[1\] VPWR VGND net3728 sg13g2_dlygate4sd3_1
X_07925_ net723 VGND VPWR net1902 i_exotiny._1924_\[18\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
Xhold49 _00078_ VPWR VGND net1876 sg13g2_dlygate4sd3_1
Xhold1945 i_exotiny.gpo\[0\] VPWR VGND net3772 sg13g2_dlygate4sd3_1
Xhold1912 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[0\]
+ VPWR VGND net3739 sg13g2_dlygate4sd3_1
Xhold1934 i_exotiny._0550_ VPWR VGND net3761 sg13g2_dlygate4sd3_1
Xhold1923 i_exotiny._1611_\[25\] VPWR VGND net3750 sg13g2_dlygate4sd3_1
Xhold1978 i_exotiny.i_wb_spi.sck_r VPWR VGND net3805 sg13g2_dlygate4sd3_1
Xhold1956 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[4\] VPWR VGND net3783
+ sg13g2_dlygate4sd3_1
Xhold1967 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[3\] VPWR VGND net3794
+ sg13g2_dlygate4sd3_1
X_07856_ net2273 net879 _03222_ _03226_ VPWR VGND sg13g2_mux2_1
X_06807_ net2012 net1096 _02827_ VPWR VGND sg13g2_nor2_1
XFILLER_25_810 VPWR VGND sg13g2_fill_2
X_07787_ i_exotiny._0023_\[1\] net3203 net895 _01266_ VPWR VGND sg13g2_mux2_1
X_04999_ _01392_ net1180 _01731_ VPWR VGND sg13g2_nor2_1
Xhold1989 i_exotiny._1618_\[3\] VPWR VGND net3816 sg13g2_dlygate4sd3_1
X_06738_ VGND VPWR _01410_ net1190 _02768_ net1169 sg13g2_a21oi_1
X_08875__1107 VPWR VGND net1527 sg13g2_tiehi
XFILLER_43_117 VPWR VGND sg13g2_fill_1
X_08911__1071 VPWR VGND net1491 sg13g2_tiehi
X_08408_ net277 VGND VPWR net2270 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[7\]
+ clknet_leaf_97_clk_regs sg13g2_dfrbpq_1
X_09217__762 VPWR VGND net762 sg13g2_tiehi
X_06669_ _02688_ VPWR _02707_ VGND _02465_ _02470_ sg13g2_o21ai_1
X_08339_ net339 VGND VPWR _00420_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[9\]
+ clknet_leaf_95_clk_regs sg13g2_dfrbpq_1
X_08578__1406 VPWR VGND net1826 sg13g2_tiehi
X_09148__834 VPWR VGND net834 sg13g2_tiehi
XFILLER_106_664 VPWR VGND sg13g2_decap_8
XFILLER_105_130 VPWR VGND sg13g2_decap_8
Xfanout1003 net1004 net1003 VPWR VGND sg13g2_buf_8
Xclkbuf_regs_0_clk clk clk_regs VPWR VGND sg13g2_buf_8
XFILLER_0_931 VPWR VGND sg13g2_decap_8
Xfanout1014 net1016 net1014 VPWR VGND sg13g2_buf_8
Xfanout1025 net1027 net1025 VPWR VGND sg13g2_buf_8
Xfanout1036 net1037 net1036 VPWR VGND sg13g2_buf_8
X_09224__755 VPWR VGND net755 sg13g2_tiehi
Xfanout1047 _02527_ net1047 VPWR VGND sg13g2_buf_8
XFILLER_102_881 VPWR VGND sg13g2_decap_8
Xfanout1058 net1059 net1058 VPWR VGND sg13g2_buf_2
XFILLER_59_250 VPWR VGND sg13g2_fill_2
Xfanout1069 net1070 net1069 VPWR VGND sg13g2_buf_8
XFILLER_101_380 VPWR VGND sg13g2_decap_8
XFILLER_48_957 VPWR VGND sg13g2_fill_2
XFILLER_19_82 VPWR VGND sg13g2_fill_2
XFILLER_90_713 VPWR VGND sg13g2_fill_1
X_08448__232 VPWR VGND net232 sg13g2_tiehi
XFILLER_27_180 VPWR VGND sg13g2_fill_1
XFILLER_34_117 VPWR VGND sg13g2_fill_2
X_09155__827 VPWR VGND net827 sg13g2_tiehi
XFILLER_35_92 VPWR VGND sg13g2_fill_2
X_09231__748 VPWR VGND net748 sg13g2_tiehi
X_08731__1257 VPWR VGND net1677 sg13g2_tiehi
Xhold508 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[12\]
+ VPWR VGND net2335 sg13g2_dlygate4sd3_1
Xhold519 _01284_ VPWR VGND net2346 sg13g2_dlygate4sd3_1
X_08455__225 VPWR VGND net225 sg13g2_tiehi
XFILLER_98_846 VPWR VGND sg13g2_decap_8
X_08953__1029 VPWR VGND net1449 sg13g2_tiehi
Xclkbuf_leaf_147_clk_regs clknet_5_16__leaf_clk_regs clknet_leaf_147_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_97_345 VPWR VGND sg13g2_decap_8
Xhold1219 _00813_ VPWR VGND net3046 sg13g2_dlygate4sd3_1
X_05971_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[1\] _02474_ _02492_
+ VPWR VGND net1262 sg13g2_nand3b_1
X_07710_ net3176 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[7\]
+ net995 _01206_ VPWR VGND sg13g2_mux2_1
Xhold1208 _00773_ VPWR VGND net3035 sg13g2_dlygate4sd3_1
X_08690_ net1718 VGND VPWR net1995 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[17\]
+ clknet_leaf_121_clk_regs sg13g2_dfrbpq_1
X_04922_ _01614_ _01620_ _01654_ VPWR VGND sg13g2_nor2_2
XFILLER_93_584 VPWR VGND sg13g2_fill_1
XFILLER_65_253 VPWR VGND sg13g2_fill_1
X_04853_ VGND VPWR net1072 _01588_ i_exotiny._1902_\[3\] _01589_ sg13g2_a21oi_1
X_07641_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[14\]
+ net3338 net897 _01149_ VPWR VGND sg13g2_mux2_1
X_07572_ net3201 net1830 _03153_ VPWR VGND sg13g2_nor2_1
X_08462__218 VPWR VGND net218 sg13g2_tiehi
X_06523_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[12\]
+ net2874 net933 _00598_ VPWR VGND sg13g2_mux2_1
X_04784_ VPWR VGND _01533_ net1273 _01437_ net1224 _01534_ net1234 sg13g2_a221oi_1
XFILLER_90_1028 VPWR VGND sg13g2_fill_1
XFILLER_90_1017 VPWR VGND sg13g2_decap_8
X_06454_ net3166 net2679 net935 _00541_ VPWR VGND sg13g2_mux2_1
X_09242_ net565 VGND VPWR net2135 i_exotiny._0022_\[0\] clknet_leaf_126_clk_regs sg13g2_dfrbpq_2
X_08707__1281 VPWR VGND net1701 sg13g2_tiehi
X_05405_ VGND VPWR i_exotiny._2034_\[5\] _02115_ _02118_ i_exotiny._2034_\[6\] sg13g2_a21oi_1
X_09173_ net809 VGND VPWR _01228_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[29\]
+ clknet_leaf_171_clk_regs sg13g2_dfrbpq_1
X_06385_ net3775 _01484_ _01489_ _01521_ _02574_ VPWR VGND sg13g2_nor4_1
X_08182__495 VPWR VGND net495 sg13g2_tiehi
X_05336_ _02060_ _02041_ _02047_ _01979_ _01978_ VPWR VGND sg13g2_a22oi_1
X_08124_ net570 VGND VPWR _00205_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[29\]
+ clknet_leaf_122_clk_regs sg13g2_dfrbpq_1
X_08055_ net639 VGND VPWR _00136_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[24\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
X_08602__1374 VPWR VGND net1794 sg13g2_tiehi
X_05267_ _01993_ _01787_ i_exotiny._0031_\[0\] _01779_ i_exotiny._0020_\[0\] VPWR
+ VGND sg13g2_a22oi_1
Xoutput39 net39 uo_out[5] VPWR VGND sg13g2_buf_1
Xoutput28 net28 uio_out[2] VPWR VGND sg13g2_buf_1
X_05198_ _01926_ _01782_ i_exotiny._0037_\[1\] _01763_ i_exotiny._0029_\[1\] VPWR
+ VGND sg13g2_a22oi_1
X_07006_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[10\]
+ net3034 net921 _00773_ VPWR VGND sg13g2_mux2_1
XFILLER_89_835 VPWR VGND sg13g2_fill_2
X_08929__1053 VPWR VGND net1473 sg13g2_tiehi
X_08957_ net1445 VGND VPWR net3472 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[23\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
Xhold1720 i_exotiny._0315_\[14\] VPWR VGND net3547 sg13g2_dlygate4sd3_1
Xhold1742 i_exotiny.i_wdg_top.clk_div_inst.cnt\[18\] VPWR VGND net3569 sg13g2_dlygate4sd3_1
X_07908_ net1175 VGND VPWR net1127 i_exotiny._3871_ clknet_leaf_35_clk_regs sg13g2_dfrbpq_2
X_08888_ net1514 VGND VPWR net1938 i_exotiny.i_wb_spi.dat_rx_r\[18\] clknet_leaf_62_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_29_434 VPWR VGND sg13g2_fill_1
Xhold1731 i_exotiny._1160_\[17\] VPWR VGND net3558 sg13g2_dlygate4sd3_1
Xhold1753 i_exotiny._0079_\[4\] VPWR VGND net3580 sg13g2_dlygate4sd3_1
XFILLER_57_765 VPWR VGND sg13g2_fill_1
Xhold1764 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[0\] VPWR VGND net3591
+ sg13g2_dlygate4sd3_1
Xhold1775 i_exotiny._1611_\[9\] VPWR VGND net3602 sg13g2_dlygate4sd3_1
Xhold1786 _01085_ VPWR VGND net3613 sg13g2_dlygate4sd3_1
X_07839_ net3446 net3222 net983 _01312_ VPWR VGND sg13g2_mux2_1
Xhold1797 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data[0]
+ VPWR VGND net3624 sg13g2_dlygate4sd3_1
XFILLER_9_806 VPWR VGND sg13g2_fill_1
XFILLER_106_461 VPWR VGND sg13g2_decap_8
XFILLER_97_65 VPWR VGND sg13g2_fill_2
XFILLER_79_334 VPWR VGND sg13g2_fill_2
X_08749__1239 VPWR VGND net1659 sg13g2_tiehi
XFILLER_95_849 VPWR VGND sg13g2_decap_8
XFILLER_94_326 VPWR VGND sg13g2_decap_8
XFILLER_94_359 VPWR VGND sg13g2_fill_2
X_09022__960 VPWR VGND net1380 sg13g2_tiehi
X_06170_ net3441 net3435 net952 _00332_ VPWR VGND sg13g2_mux2_1
Xhold305 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[26\]
+ VPWR VGND net2132 sg13g2_dlygate4sd3_1
XFILLER_7_85 VPWR VGND sg13g2_fill_1
Xhold316 _01307_ VPWR VGND net2143 sg13g2_dlygate4sd3_1
X_05121_ _01851_ _01771_ i_exotiny._0016_\[2\] _01763_ i_exotiny._0029_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold338 _00133_ VPWR VGND net2165 sg13g2_dlygate4sd3_1
Xhold327 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[12\]
+ VPWR VGND net2154 sg13g2_dlygate4sd3_1
Xhold349 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[23\]
+ VPWR VGND net2176 sg13g2_dlygate4sd3_1
X_05052_ net1238 net1241 net1235 _01784_ VGND VPWR _01759_ sg13g2_nor4_2
X_08577__49 VPWR VGND net49 sg13g2_tiehi
XFILLER_30_0 VPWR VGND sg13g2_fill_2
X_09207__772 VPWR VGND net772 sg13g2_tiehi
X_08811_ net1597 VGND VPWR _00869_ i_exotiny.i_wb_spi.state_r\[10\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
Xhold1005 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[13\]
+ VPWR VGND net2832 sg13g2_dlygate4sd3_1
Xhold1027 _01264_ VPWR VGND net2854 sg13g2_dlygate4sd3_1
X_08742_ net1666 VGND VPWR net2294 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[5\]
+ clknet_leaf_86_clk_regs sg13g2_dfrbpq_1
X_05954_ net2892 net2456 net969 _00163_ VPWR VGND sg13g2_mux2_1
Xhold1049 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[17\]
+ VPWR VGND net2876 sg13g2_dlygate4sd3_1
Xhold1016 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[10\]
+ VPWR VGND net2843 sg13g2_dlygate4sd3_1
Xhold1038 _00641_ VPWR VGND net2865 sg13g2_dlygate4sd3_1
XFILLER_94_860 VPWR VGND sg13g2_fill_2
Xclkbuf_4_7_0_clk_regs clknet_0_clk_regs clknet_4_7_0_clk_regs VPWR VGND sg13g2_buf_8
X_08673_ net1735 VGND VPWR _00731_ i_exotiny._0034_\[0\] clknet_leaf_102_clk_regs
+ sg13g2_dfrbpq_2
X_04905_ net1258 net1260 net1222 _01637_ VGND VPWR _01623_ sg13g2_nor4_2
XFILLER_38_231 VPWR VGND sg13g2_fill_2
X_07624_ VPWR _01134_ _03186_ VGND sg13g2_inv_1
X_05885_ _02465_ _02470_ _02471_ VPWR VGND sg13g2_nor2_2
XFILLER_26_437 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_44_clk_regs clknet_5_11__leaf_clk_regs clknet_leaf_44_clk_regs VPWR VGND
+ sg13g2_buf_8
X_04836_ i_exotiny.i_wb_spi.cnt_presc_r\[6\] _01575_ _01576_ VPWR VGND sg13g2_nor2_1
X_09138__844 VPWR VGND net844 sg13g2_tiehi
X_07555_ net3681 _03140_ _03142_ VPWR VGND sg13g2_and2_1
X_04767_ net1270 net1273 _01518_ VPWR VGND sg13g2_nor2_1
X_06506_ _02618_ net2341 net1025 _00584_ VPWR VGND sg13g2_mux2_1
XFILLER_22_643 VPWR VGND sg13g2_fill_2
X_07486_ net3692 net903 _03110_ VPWR VGND sg13g2_nor2_1
X_06437_ net2777 net3291 net937 _00524_ VPWR VGND sg13g2_mux2_1
X_09214__765 VPWR VGND net765 sg13g2_tiehi
X_09225_ net754 VGND VPWR _01280_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[15\]
+ clknet_leaf_134_clk_regs sg13g2_dfrbpq_1
XFILLER_21_153 VPWR VGND sg13g2_fill_1
X_04698_ _01456_ net1248 net1247 VPWR VGND sg13g2_nand2_1
X_06368_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[27\]
+ net2515 net1031 _00498_ VPWR VGND sg13g2_mux2_1
X_09156_ net826 VGND VPWR _01211_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[12\]
+ clknet_leaf_175_clk_regs sg13g2_dfrbpq_1
X_06299_ _02555_ net2424 net939 _00440_ VPWR VGND sg13g2_mux2_1
X_08107_ net587 VGND VPWR _00188_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[12\]
+ clknet_leaf_101_clk_regs sg13g2_dfrbpq_1
X_09087_ net1315 VGND VPWR net2860 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[7\]
+ clknet_leaf_145_clk_regs sg13g2_dfrbpq_1
X_05319_ VPWR VGND _02012_ net1109 _01988_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[0\]
+ _02044_ net1107 sg13g2_a221oi_1
X_08038_ net656 VGND VPWR _00119_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[7\]
+ clknet_leaf_55_clk_regs sg13g2_dfrbpq_1
Xhold850 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[5\]
+ VPWR VGND net2677 sg13g2_dlygate4sd3_1
X_09145__837 VPWR VGND net837 sg13g2_tiehi
Xhold861 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[8\]
+ VPWR VGND net2688 sg13g2_dlygate4sd3_1
Xhold872 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[22\]
+ VPWR VGND net2699 sg13g2_dlygate4sd3_1
XFILLER_104_965 VPWR VGND sg13g2_decap_8
XFILLER_89_643 VPWR VGND sg13g2_fill_2
XFILLER_88_120 VPWR VGND sg13g2_fill_1
Xhold894 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[7\]
+ VPWR VGND net2721 sg13g2_dlygate4sd3_1
Xhold883 _00306_ VPWR VGND net2710 sg13g2_dlygate4sd3_1
XFILLER_103_486 VPWR VGND sg13g2_decap_8
XFILLER_88_175 VPWR VGND sg13g2_fill_1
XFILLER_88_153 VPWR VGND sg13g2_fill_1
X_09221__758 VPWR VGND net758 sg13g2_tiehi
Xhold1550 i_exotiny._0315_\[30\] VPWR VGND net3377 sg13g2_dlygate4sd3_1
Xhold1561 i_exotiny._1611_\[11\] VPWR VGND net3388 sg13g2_dlygate4sd3_1
XFILLER_83_23 VPWR VGND sg13g2_fill_1
Xhold1572 i_exotiny.i_wb_spi.cnt_hbit_r\[2\] VPWR VGND net3399 sg13g2_dlygate4sd3_1
Xhold1594 _01316_ VPWR VGND net3421 sg13g2_dlygate4sd3_1
Xhold1583 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[7\]
+ VPWR VGND net3410 sg13g2_dlygate4sd3_1
XFILLER_17_459 VPWR VGND sg13g2_fill_2
XFILLER_5_875 VPWR VGND sg13g2_decap_8
XFILLER_4_352 VPWR VGND sg13g2_fill_2
X_08452__228 VPWR VGND net228 sg13g2_tiehi
X_08870__1112 VPWR VGND net1532 sg13g2_tiehi
X_05670_ VGND VPWR net1062 _02323_ _00043_ _02321_ sg13g2_a21oi_1
XFILLER_91_896 VPWR VGND sg13g2_fill_2
XFILLER_63_598 VPWR VGND sg13g2_fill_2
X_04621_ _01383_ net1230 VPWR VGND sg13g2_inv_2
XFILLER_17_971 VPWR VGND sg13g2_fill_2
XFILLER_16_481 VPWR VGND sg13g2_fill_1
X_07340_ _03004_ _02995_ _03000_ VPWR VGND sg13g2_nand2_2
X_07271_ net3049 net874 _02972_ _02977_ VPWR VGND sg13g2_mux2_1
X_08144__541 VPWR VGND net541 sg13g2_tiehi
X_09010_ net1392 VGND VPWR _01068_ i_exotiny._0079_\[3\] clknet_leaf_161_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_78_0 VPWR VGND sg13g2_fill_1
X_06222_ net2871 net883 _02540_ _02543_ VPWR VGND sg13g2_mux2_1
X_06153_ i_exotiny._0028_\[1\] net3393 net951 _00315_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_162_clk_regs clknet_5_6__leaf_clk_regs clknet_leaf_162_clk_regs VPWR
+ VGND sg13g2_buf_8
Xhold113 _00039_ VPWR VGND net1940 sg13g2_dlygate4sd3_1
Xhold124 i_exotiny.i_wb_spi.dat_rx_r\[16\] VPWR VGND net1951 sg13g2_dlygate4sd3_1
Xhold135 _01232_ VPWR VGND net1962 sg13g2_dlygate4sd3_1
Xhold102 _00057_ VPWR VGND net1929 sg13g2_dlygate4sd3_1
X_05104_ _01833_ _01832_ _01828_ _01834_ VPWR VGND sg13g2_a21o_2
Xhold146 _00059_ VPWR VGND net1973 sg13g2_dlygate4sd3_1
X_06084_ net2843 net3131 net958 _00260_ VPWR VGND sg13g2_mux2_1
Xhold168 _00748_ VPWR VGND net1995 sg13g2_dlygate4sd3_1
Xhold157 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[2\] VPWR
+ VGND net1984 sg13g2_dlygate4sd3_1
Xhold179 i_exotiny._1924_\[10\] VPWR VGND net2006 sg13g2_dlygate4sd3_1
X_05035_ net1239 net1240 net1220 _01767_ VGND VPWR _01754_ sg13g2_nor4_2
XFILLER_101_913 VPWR VGND sg13g2_decap_8
XFILLER_99_996 VPWR VGND sg13g2_decap_8
XFILLER_85_101 VPWR VGND sg13g2_fill_2
XFILLER_58_315 VPWR VGND sg13g2_fill_1
XFILLER_100_423 VPWR VGND sg13g2_decap_8
XFILLER_98_495 VPWR VGND sg13g2_decap_8
XFILLER_85_145 VPWR VGND sg13g2_fill_2
X_06986_ net2450 net889 _02922_ _02924_ VPWR VGND sg13g2_mux2_1
XFILLER_96_1012 VPWR VGND sg13g2_decap_8
X_05937_ i_exotiny._0020_\[2\] net2168 net966 _00146_ VPWR VGND sg13g2_mux2_1
XFILLER_2_1027 VPWR VGND sg13g2_fill_2
X_08725_ net1683 VGND VPWR net3396 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[20\]
+ clknet_leaf_119_clk_regs sg13g2_dfrbpq_1
X_05868_ _02455_ net3370 net1056 _00109_ VPWR VGND sg13g2_mux2_1
X_08544__112 VPWR VGND net112 sg13g2_tiehi
X_08656_ net1741 VGND VPWR _00724_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[25\]
+ clknet_leaf_148_clk_regs sg13g2_dfrbpq_1
X_07607_ net1205 net3236 _03175_ _01128_ VPWR VGND sg13g2_nor3_1
X_04819_ net22 _01557_ _01559_ VPWR VGND sg13g2_nand2_2
X_08587_ net1810 VGND VPWR i_exotiny._1265_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_hlt_pc_ccx
+ clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
X_05799_ VPWR VGND _01605_ _01421_ _01533_ _01431_ _02416_ _01433_ sg13g2_a221oi_1
X_07538_ _03131_ _01362_ _01442_ VPWR VGND sg13g2_nand2_1
X_07469_ _03101_ _03102_ _03078_ _01063_ VPWR VGND sg13g2_nand3_1
X_09208_ net771 VGND VPWR _01263_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[30\]
+ clknet_leaf_76_clk_regs sg13g2_dfrbpq_1
XFILLER_6_639 VPWR VGND sg13g2_decap_4
X_09139_ net843 VGND VPWR net2210 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[27\]
+ clknet_leaf_156_clk_regs sg13g2_dfrbpq_1
X_09012__970 VPWR VGND net1390 sg13g2_tiehi
X_08551__105 VPWR VGND net105 sg13g2_tiehi
XFILLER_89_440 VPWR VGND sg13g2_fill_2
Xhold680 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[16\]
+ VPWR VGND net2507 sg13g2_dlygate4sd3_1
XFILLER_2_845 VPWR VGND sg13g2_decap_8
XFILLER_104_762 VPWR VGND sg13g2_decap_8
Xhold691 _01225_ VPWR VGND net2518 sg13g2_dlygate4sd3_1
XFILLER_103_283 VPWR VGND sg13g2_decap_8
XFILLER_45_510 VPWR VGND sg13g2_fill_1
Xhold1380 _00437_ VPWR VGND net3207 sg13g2_dlygate4sd3_1
Xhold1391 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[18\]
+ VPWR VGND net3218 sg13g2_dlygate4sd3_1
XFILLER_72_395 VPWR VGND sg13g2_fill_1
X_08699__1289 VPWR VGND net1709 sg13g2_tiehi
XFILLER_14_974 VPWR VGND sg13g2_decap_8
XFILLER_43_81 VPWR VGND sg13g2_fill_2
Xclkbuf_5_22__f_clk_regs clknet_4_11_0_clk_regs clknet_5_22__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_10678_ net1827 net29 VPWR VGND sg13g2_buf_1
XFILLER_99_226 VPWR VGND sg13g2_decap_8
XFILLER_99_248 VPWR VGND sg13g2_decap_8
X_09128__854 VPWR VGND net854 sg13g2_tiehi
XFILLER_96_900 VPWR VGND sg13g2_decap_8
X_06840_ net1170 VPWR _02854_ VGND net3638 net1185 sg13g2_o21ai_1
XFILLER_96_977 VPWR VGND sg13g2_decap_8
X_06771_ _02795_ VPWR _02796_ VGND net3759 net1190 sg13g2_o21ai_1
XFILLER_36_521 VPWR VGND sg13g2_fill_2
X_08510_ net170 VGND VPWR net2342 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[30\]
+ clknet_leaf_71_clk_regs sg13g2_dfrbpq_1
X_05722_ VGND VPWR net1058 _02362_ _00056_ _02360_ sg13g2_a21oi_1
X_05653_ VGND VPWR i_exotiny._1614_\[1\] net1125 _02311_ _02310_ sg13g2_a21oi_1
X_08441_ net244 VGND VPWR _00515_ i_exotiny._2025_\[3\] clknet_leaf_30_clk_regs sg13g2_dfrbpq_2
XFILLER_90_181 VPWR VGND sg13g2_fill_1
X_04604_ net3624 _01366_ VPWR VGND sg13g2_inv_4
X_08372_ net306 VGND VPWR _00453_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[10\]
+ clknet_leaf_137_clk_regs sg13g2_dfrbpq_1
X_05584_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[0\].i_hadd.a_i
+ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r[0] i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[1\].i_hadd.a_i
+ _02259_ VPWR VGND sg13g2_nand3_1
X_09135__847 VPWR VGND net847 sg13g2_tiehi
XFILLER_32_771 VPWR VGND sg13g2_fill_2
X_07323_ net3761 net3457 net1151 _01032_ VPWR VGND sg13g2_mux2_1
X_07254_ net2713 net2924 net1005 _00977_ VPWR VGND sg13g2_mux2_1
X_06205_ net2643 net3186 net946 _00360_ VPWR VGND sg13g2_mux2_1
X_09211__768 VPWR VGND net768 sg13g2_tiehi
X_07185_ net1281 VPWR _02957_ VGND net3772 _02956_ sg13g2_o21ai_1
XFILLER_105_515 VPWR VGND sg13g2_decap_8
X_08744__1244 VPWR VGND net1664 sg13g2_tiehi
XFILLER_2_119 VPWR VGND sg13g2_fill_1
X_06136_ net2333 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[23\]
+ net1044 _00305_ VPWR VGND sg13g2_mux2_1
X_06067_ _02515_ net2800 net963 _00248_ VPWR VGND sg13g2_mux2_1
XFILLER_99_782 VPWR VGND sg13g2_fill_2
XFILLER_87_900 VPWR VGND sg13g2_fill_1
X_05018_ _01602_ VPWR _01750_ VGND net1174 _01499_ sg13g2_o21ai_1
XFILLER_98_292 VPWR VGND sg13g2_decap_8
XFILLER_100_220 VPWR VGND sg13g2_decap_8
XFILLER_87_999 VPWR VGND sg13g2_decap_8
XFILLER_74_616 VPWR VGND sg13g2_fill_1
XFILLER_86_487 VPWR VGND sg13g2_fill_2
XFILLER_74_627 VPWR VGND sg13g2_fill_2
XFILLER_58_189 VPWR VGND sg13g2_decap_4
X_06969_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[11\]
+ net3288 net1020 _00742_ VPWR VGND sg13g2_mux2_1
XFILLER_100_297 VPWR VGND sg13g2_decap_8
XFILLER_73_159 VPWR VGND sg13g2_fill_1
X_08708_ net1700 VGND VPWR net2094 i_exotiny._0032_\[3\] clknet_leaf_117_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_55_896 VPWR VGND sg13g2_fill_2
XFILLER_54_373 VPWR VGND sg13g2_decap_8
X_08966__1016 VPWR VGND net1436 sg13g2_tiehi
X_08639_ net1758 VGND VPWR net2689 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[8\]
+ clknet_leaf_143_clk_regs sg13g2_dfrbpq_1
XFILLER_42_557 VPWR VGND sg13g2_decap_4
XFILLER_70_1026 VPWR VGND sg13g2_fill_2
XFILLER_7_926 VPWR VGND sg13g2_decap_8
XFILLER_11_988 VPWR VGND sg13g2_decap_8
X_07980__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_8_0 VPWR VGND sg13g2_fill_2
XFILLER_104_570 VPWR VGND sg13g2_fill_1
XFILLER_77_421 VPWR VGND sg13g2_fill_1
XFILLER_93_914 VPWR VGND sg13g2_decap_8
X_08615__1361 VPWR VGND net1781 sg13g2_tiehi
Xfanout990 net992 net990 VPWR VGND sg13g2_buf_8
XFILLER_65_649 VPWR VGND sg13g2_fill_1
Xclkbuf_5_6__f_clk_regs clknet_4_3_0_clk_regs clknet_5_6__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_45_362 VPWR VGND sg13g2_fill_1
X_08822__1166 VPWR VGND net1586 sg13g2_tiehi
XFILLER_20_207 VPWR VGND sg13g2_fill_2
XFILLER_86_1011 VPWR VGND sg13g2_decap_8
X_08395__535 VPWR VGND net535 sg13g2_tiehi
Xclkload22 clkload22/Y clknet_leaf_27_clk_regs VPWR VGND sg13g2_inv_2
X_08141__544 VPWR VGND net544 sg13g2_tiehi
Xclkload33 VPWR clkload33/Y clknet_leaf_156_clk_regs VGND sg13g2_inv_1
Xclkload11 clknet_leaf_10_clk_regs clkload11/Y VPWR VGND sg13g2_inv_4
XFILLER_102_518 VPWR VGND sg13g2_decap_8
X_08990_ net1412 VGND VPWR net3527 i_exotiny._1160_\[11\] clknet_leaf_161_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_102_529 VPWR VGND sg13g2_fill_1
X_07941_ net85 VGND VPWR _00006_ i_exotiny._1793_ clknet_leaf_27_clk_regs sg13g2_dfrbpq_2
XFILLER_96_763 VPWR VGND sg13g2_fill_2
X_07872_ net3268 net3445 net981 _01339_ VPWR VGND sg13g2_mux2_1
X_06823_ net1132 _02838_ _02839_ _02840_ VPWR VGND sg13g2_nor3_1
X_06754_ _02782_ _02719_ net3559 net1068 net3142 VPWR VGND sg13g2_a22oi_1
X_05705_ net1924 net1058 _02350_ VPWR VGND sg13g2_nor2_1
XFILLER_93_1026 VPWR VGND sg13g2_fill_2
XFILLER_92_991 VPWR VGND sg13g2_decap_8
XFILLER_63_170 VPWR VGND sg13g2_fill_1
X_06685_ i_exotiny._0315_\[3\] net1233 _01391_ _02722_ VPWR VGND sg13g2_nor3_1
X_09002__980 VPWR VGND net1400 sg13g2_tiehi
X_05636_ net1119 net1943 _02298_ VPWR VGND sg13g2_nor2b_1
X_08424_ net261 VGND VPWR net2516 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[23\]
+ clknet_leaf_96_clk_regs sg13g2_dfrbpq_1
X_08355_ net323 VGND VPWR _00436_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[25\]
+ clknet_leaf_94_clk_regs sg13g2_dfrbpq_1
X_05567_ VGND VPWR net3523 net3677 _02248_ _02247_ sg13g2_a21oi_1
Xclkload5 clknet_5_27__leaf_clk_regs clkload5/X VPWR VGND sg13g2_buf_8
X_07306_ net2880 _02981_ net908 _01021_ VPWR VGND sg13g2_mux2_1
X_08286_ net392 VGND VPWR net2376 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[20\]
+ clknet_leaf_100_clk_regs sg13g2_dfrbpq_1
XFILLER_50_16 VPWR VGND sg13g2_decap_8
X_05498_ _02191_ VPWR i_exotiny._1611_\[13\] VGND net1076 _02193_ sg13g2_o21ai_1
X_07237_ net3314 net3341 net1004 _00960_ VPWR VGND sg13g2_mux2_1
X_07168_ net2660 net3160 net1008 _00916_ VPWR VGND sg13g2_mux2_1
XFILLER_4_918 VPWR VGND sg13g2_decap_8
XFILLER_106_846 VPWR VGND sg13g2_decap_8
XFILLER_105_312 VPWR VGND sg13g2_decap_8
X_06119_ net2691 net2961 net1047 _00288_ VPWR VGND sg13g2_mux2_1
XFILLER_1_7 VPWR VGND sg13g2_decap_8
X_07099_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[27\]
+ net2216 net914 _00854_ VPWR VGND sg13g2_mux2_1
XFILLER_105_389 VPWR VGND sg13g2_decap_8
Xfanout1229 i_exotiny.i_wdg_top.clk_div_inst.cnt\[19\] net1229 VPWR VGND sg13g2_buf_1
XFILLER_8_1000 VPWR VGND sg13g2_decap_8
Xfanout1207 net1209 net1207 VPWR VGND sg13g2_buf_8
Xfanout1218 _01489_ net1218 VPWR VGND sg13g2_buf_8
XFILLER_101_584 VPWR VGND sg13g2_fill_2
XFILLER_43_811 VPWR VGND sg13g2_fill_2
XFILLER_42_332 VPWR VGND sg13g2_fill_1
XFILLER_30_538 VPWR VGND sg13g2_decap_4
X_09118__864 VPWR VGND net864 sg13g2_tiehi
XFILLER_24_83 VPWR VGND sg13g2_fill_1
XFILLER_11_774 VPWR VGND sg13g2_fill_2
XFILLER_97_516 VPWR VGND sg13g2_decap_8
XFILLER_3_984 VPWR VGND sg13g2_decap_8
X_09125__857 VPWR VGND net857 sg13g2_tiehi
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_92_298 VPWR VGND sg13g2_decap_8
X_09171__811 VPWR VGND net811 sg13g2_tiehi
X_06470_ _02613_ net3346 net935 _00553_ VPWR VGND sg13g2_mux2_1
XFILLER_33_387 VPWR VGND sg13g2_fill_2
X_05421_ VGND VPWR _01387_ net1234 _02130_ net1244 sg13g2_a21oi_1
X_08140_ net545 VGND VPWR _00221_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[4\]
+ clknet_leaf_131_clk_regs sg13g2_dfrbpq_1
X_05352_ _02074_ net1263 _01402_ VPWR VGND sg13g2_nand2_1
X_08071_ net623 VGND VPWR _00152_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[8\]
+ clknet_leaf_89_clk_regs sg13g2_dfrbpq_1
X_05283_ VPWR VGND i_exotiny._0037_\[0\] _02008_ _01782_ i_exotiny._0032_\[0\] _02009_
+ _01767_ sg13g2_a221oi_1
Xclkbuf_leaf_69_clk_regs clknet_5_25__leaf_clk_regs clknet_leaf_69_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07022_ net2111 net3077 net920 _00789_ VPWR VGND sg13g2_mux2_1
XFILLER_102_315 VPWR VGND sg13g2_decap_8
X_08973_ net1429 VGND VPWR _01031_ i_exotiny._0571_ clknet_leaf_12_clk_regs sg13g2_dfrbpq_2
Xhold17 i_exotiny.i_wb_spi.state_r\[29\] VPWR VGND net1844 sg13g2_dlygate4sd3_1
Xhold28 i_exotiny.i_wb_spi.state_r\[6\] VPWR VGND net1855 sg13g2_dlygate4sd3_1
X_07924_ net724 VGND VPWR net2032 i_exotiny._1924_\[17\] clknet_leaf_34_clk_regs sg13g2_dfrbpq_1
Xhold1902 i_exotiny._0369_\[3\] VPWR VGND net3729 sg13g2_dlygate4sd3_1
Xhold39 i_exotiny.i_wb_spi.state_r\[28\] VPWR VGND net1866 sg13g2_dlygate4sd3_1
Xhold1924 i_exotiny.i_wdg_top.o_wb_dat\[6\] VPWR VGND net3751 sg13g2_dlygate4sd3_1
Xhold1935 i_exotiny._0315_\[3\] VPWR VGND net3762 sg13g2_dlygate4sd3_1
Xhold1913 _01033_ VPWR VGND net3740 sg13g2_dlygate4sd3_1
Xhold1968 i_exotiny.i_wdg_top.o_wb_dat\[5\] VPWR VGND net3795 sg13g2_dlygate4sd3_1
Xhold1946 _02957_ VPWR VGND net3773 sg13g2_dlygate4sd3_1
X_08694__1294 VPWR VGND net1714 sg13g2_tiehi
X_07855_ _03225_ net2910 net985 _01326_ VPWR VGND sg13g2_mux2_1
Xhold1957 i_exotiny._0315_\[5\] VPWR VGND net3784 sg13g2_dlygate4sd3_1
Xhold1979 _01231_ VPWR VGND net3806 sg13g2_dlygate4sd3_1
X_06806_ VGND VPWR net3697 net1130 _02826_ _02825_ sg13g2_a21oi_1
X_07786_ i_exotiny._0023_\[0\] net3227 net894 _01265_ VPWR VGND sg13g2_mux2_1
X_04998_ _01727_ _01728_ _01709_ _01730_ VPWR VGND sg13g2_nand3_1
XFILLER_83_287 VPWR VGND sg13g2_fill_2
X_06737_ _02767_ net3714 net1183 VPWR VGND sg13g2_nand2_1
XFILLER_101_33 VPWR VGND sg13g2_fill_2
X_06668_ VPWR VGND _02706_ net1196 _02705_ _01370_ _00658_ net1154 sg13g2_a221oi_1
X_08407_ net278 VGND VPWR net3374 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[6\]
+ clknet_leaf_97_clk_regs sg13g2_dfrbpq_1
X_05619_ net1987 net1065 _02285_ VPWR VGND sg13g2_nor2_1
X_06599_ net3447 net1153 _02656_ VPWR VGND sg13g2_nor2_1
X_08338_ net340 VGND VPWR _00419_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[8\]
+ clknet_leaf_98_clk_regs sg13g2_dfrbpq_1
X_08269_ net409 VGND VPWR _00350_ i_exotiny._0033_\[3\] clknet_leaf_103_clk_regs sg13g2_dfrbpq_2
XFILLER_20_593 VPWR VGND sg13g2_fill_1
XFILLER_106_643 VPWR VGND sg13g2_decap_8
XFILLER_105_186 VPWR VGND sg13g2_decap_8
Xfanout1004 net1007 net1004 VPWR VGND sg13g2_buf_8
XFILLER_0_910 VPWR VGND sg13g2_decap_8
Xfanout1015 net1016 net1015 VPWR VGND sg13g2_buf_8
Xfanout1026 net1027 net1026 VPWR VGND sg13g2_buf_8
Xfanout1037 _02559_ net1037 VPWR VGND sg13g2_buf_8
XFILLER_102_860 VPWR VGND sg13g2_decap_8
Xfanout1059 net1060 net1059 VPWR VGND sg13g2_buf_1
XFILLER_0_987 VPWR VGND sg13g2_decap_8
Xfanout1048 net1049 net1048 VPWR VGND sg13g2_buf_8
XFILLER_71_972 VPWR VGND sg13g2_fill_2
XFILLER_43_674 VPWR VGND sg13g2_fill_1
Xhold509 _01207_ VPWR VGND net2336 sg13g2_dlygate4sd3_1
XFILLER_83_1014 VPWR VGND sg13g2_decap_8
XFILLER_97_324 VPWR VGND sg13g2_decap_8
XFILLER_3_781 VPWR VGND sg13g2_decap_8
X_08961__1021 VPWR VGND net1441 sg13g2_tiehi
X_05970_ net2505 _02491_ net966 _00175_ VPWR VGND sg13g2_mux2_1
XFILLER_32_4 VPWR VGND sg13g2_decap_4
XFILLER_100_819 VPWR VGND sg13g2_decap_8
Xhold1209 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[22\]
+ VPWR VGND net3036 sg13g2_dlygate4sd3_1
X_04921_ net1258 net1260 net1255 _01653_ VGND VPWR _01623_ sg13g2_nor4_2
XFILLER_18_2 VPWR VGND sg13g2_fill_1
X_04852_ VGND VPWR net3551 _01570_ _01589_ net1072 sg13g2_a21oi_1
Xclkbuf_leaf_116_clk_regs clknet_5_19__leaf_clk_regs clknet_leaf_116_clk_regs VPWR
+ VGND sg13g2_buf_8
X_07640_ net3190 net3311 net898 _01148_ VPWR VGND sg13g2_mux2_1
X_07571_ net1830 net1204 _01115_ VPWR VGND sg13g2_nor2_1
X_04783_ VGND VPWR _01533_ net1244 net1246 sg13g2_or2_1
X_06522_ net2590 net2606 net930 _00597_ VPWR VGND sg13g2_mux2_1
X_06453_ net2667 net2648 net938 _00540_ VPWR VGND sg13g2_mux2_1
X_09241_ net566 VGND VPWR _01296_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[31\]
+ clknet_leaf_133_clk_regs sg13g2_dfrbpq_1
X_05404_ net1112 _02117_ i_exotiny._2043_\[5\] VPWR VGND sg13g2_nor2_1
X_09172_ net810 VGND VPWR _01227_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[28\]
+ clknet_leaf_174_clk_regs sg13g2_dfrbpq_1
X_06384_ _00507_ _02572_ _02573_ VPWR VGND sg13g2_nand2_1
X_08123_ net571 VGND VPWR net3514 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[28\]
+ clknet_leaf_124_clk_regs sg13g2_dfrbpq_1
X_05335_ VGND VPWR _01976_ _01977_ _02059_ _01973_ sg13g2_a21oi_1
X_08054_ net640 VGND VPWR _00135_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[23\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
X_05266_ _01992_ _01781_ i_exotiny._0028_\[0\] _01766_ i_exotiny._0030_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_07005_ net2089 net3028 net920 _00772_ VPWR VGND sg13g2_mux2_1
Xoutput29 net29 uio_out[3] VPWR VGND sg13g2_buf_1
X_05197_ _01925_ _01786_ i_exotiny._0017_\[1\] _01769_ i_exotiny._0022_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xoutput18 net18 uio_oe[0] VPWR VGND sg13g2_buf_1
XFILLER_103_624 VPWR VGND sg13g2_fill_1
XFILLER_103_657 VPWR VGND sg13g2_decap_4
XFILLER_102_134 VPWR VGND sg13g2_fill_1
X_08956_ net1446 VGND VPWR _01014_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[22\]
+ clknet_leaf_54_clk_regs sg13g2_dfrbpq_1
X_08781__1207 VPWR VGND net1627 sg13g2_tiehi
X_09108__874 VPWR VGND net1294 sg13g2_tiehi
Xhold1710 i_exotiny._0315_\[10\] VPWR VGND net3537 sg13g2_dlygate4sd3_1
XFILLER_102_189 VPWR VGND sg13g2_decap_8
XFILLER_99_1010 VPWR VGND sg13g2_decap_8
XFILLER_97_891 VPWR VGND sg13g2_decap_8
X_07907_ net1176 VGND VPWR net3512 _00014_ clknet_leaf_37_clk_regs sg13g2_dfrbpq_1
Xhold1732 i_exotiny._1615_\[1\] VPWR VGND net3559 sg13g2_dlygate4sd3_1
X_08887_ net1515 VGND VPWR net1952 i_exotiny.i_wb_spi.dat_rx_r\[17\] clknet_leaf_59_clk_regs
+ sg13g2_dfrbpq_1
Xhold1743 i_exotiny._0315_\[29\] VPWR VGND net3570 sg13g2_dlygate4sd3_1
Xhold1721 _01084_ VPWR VGND net3548 sg13g2_dlygate4sd3_1
XFILLER_84_574 VPWR VGND sg13g2_fill_2
Xhold1787 i_exotiny._1616_\[2\] VPWR VGND net3614 sg13g2_dlygate4sd3_1
Xhold1765 _00618_ VPWR VGND net3592 sg13g2_dlygate4sd3_1
Xhold1776 i_exotiny._0314_\[5\] VPWR VGND net3603 sg13g2_dlygate4sd3_1
X_07838_ net2922 net2142 net984 _01311_ VPWR VGND sg13g2_mux2_1
Xhold1754 _01069_ VPWR VGND net3581 sg13g2_dlygate4sd3_1
Xhold1798 i_exotiny._0315_\[19\] VPWR VGND net3625 sg13g2_dlygate4sd3_1
X_07769_ net2696 net2951 net991 _01254_ VPWR VGND sg13g2_mux2_1
XFILLER_72_58 VPWR VGND sg13g2_fill_1
X_08839__1147 VPWR VGND net1567 sg13g2_tiehi
X_09115__867 VPWR VGND net867 sg13g2_tiehi
XFILLER_40_688 VPWR VGND sg13g2_decap_4
X_08554__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_106_440 VPWR VGND sg13g2_decap_8
X_09161__821 VPWR VGND net821 sg13g2_tiehi
XFILLER_94_305 VPWR VGND sg13g2_decap_8
XFILLER_48_711 VPWR VGND sg13g2_fill_1
XFILLER_48_700 VPWR VGND sg13g2_decap_8
X_08757__1231 VPWR VGND net1651 sg13g2_tiehi
XFILLER_0_784 VPWR VGND sg13g2_decap_8
X_08979__1003 VPWR VGND net1423 sg13g2_tiehi
X_05120_ _01850_ _01784_ i_exotiny._0042_\[2\] _01769_ i_exotiny._0022_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold306 _01255_ VPWR VGND net2133 sg13g2_dlygate4sd3_1
XFILLER_7_383 VPWR VGND sg13g2_fill_2
Xhold317 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[13\]
+ VPWR VGND net2144 sg13g2_dlygate4sd3_1
Xhold339 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[6\]
+ VPWR VGND net2166 sg13g2_dlygate4sd3_1
Xhold328 _00184_ VPWR VGND net2155 sg13g2_dlygate4sd3_1
X_05051_ i_exotiny._0079_\[2\] i_exotiny._0079_\[3\] net1235 _01783_ VGND VPWR _01762_
+ sg13g2_nor4_2
XFILLER_97_132 VPWR VGND sg13g2_fill_2
X_08810_ net1598 VGND VPWR _00868_ i_exotiny.i_wb_spi.state_r\[9\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_100_627 VPWR VGND sg13g2_fill_2
Xhold1006 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[9\]
+ VPWR VGND net2833 sg13g2_dlygate4sd3_1
XFILLER_23_0 VPWR VGND sg13g2_fill_1
X_08741_ net1667 VGND VPWR _00799_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[4\]
+ clknet_leaf_80_clk_regs sg13g2_dfrbpq_1
X_05953_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[18\]
+ net2406 net967 _00162_ VPWR VGND sg13g2_mux2_1
Xhold1039 i_exotiny._0017_\[2\] VPWR VGND net2866 sg13g2_dlygate4sd3_1
Xhold1028 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[23\]
+ VPWR VGND net2855 sg13g2_dlygate4sd3_1
Xhold1017 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[16\]
+ VPWR VGND net2844 sg13g2_dlygate4sd3_1
X_08672_ net1203 VGND VPWR i_exotiny._2043_\[9\] i_exotiny._2034_\[9\] net1229 sg13g2_dfrbpq_2
X_04904_ net1258 net1260 _01614_ _01636_ VPWR VGND sg13g2_nor3_2
X_05884_ VPWR VGND _02428_ net1184 _02469_ _02466_ _02470_ _02467_ sg13g2_a221oi_1
X_07623_ _03185_ VPWR _03186_ VGND net1228 _03183_ sg13g2_o21ai_1
XFILLER_38_287 VPWR VGND sg13g2_fill_1
XFILLER_81_555 VPWR VGND sg13g2_fill_2
XFILLER_81_533 VPWR VGND sg13g2_fill_2
X_04835_ _01575_ _01574_ i_exotiny.i_wb_spi.cnt_presc_r\[5\] VPWR VGND sg13g2_nand2b_1
X_07554_ _03140_ _03141_ _01109_ VPWR VGND sg13g2_nor2_1
X_04766_ VGND VPWR _01517_ net1181 net1219 sg13g2_or2_1
XFILLER_41_408 VPWR VGND sg13g2_fill_2
X_06505_ i_exotiny._0041_\[2\] net878 _02614_ _02618_ VPWR VGND sg13g2_mux2_1
X_04697_ _01446_ VPWR _01455_ VGND net1266 _01454_ sg13g2_o21ai_1
X_07485_ _03109_ VPWR _01072_ VGND _01386_ net906 sg13g2_o21ai_1
Xclkbuf_leaf_84_clk_regs clknet_5_30__leaf_clk_regs clknet_leaf_84_clk_regs VPWR VGND
+ sg13g2_buf_8
X_09224_ net755 VGND VPWR net2752 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[14\]
+ clknet_leaf_136_clk_regs sg13g2_dfrbpq_1
X_06436_ net3037 net3064 net936 _00523_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_13_clk_regs clknet_5_3__leaf_clk_regs clknet_leaf_13_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06367_ net2196 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[22\]
+ net1031 _00497_ VPWR VGND sg13g2_mux2_1
X_09155_ net827 VGND VPWR _01210_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[11\]
+ clknet_leaf_173_clk_regs sg13g2_dfrbpq_1
X_06298_ i_exotiny._0016_\[1\] net884 _02552_ _02555_ VPWR VGND sg13g2_mux2_1
X_08835__1153 VPWR VGND net1573 sg13g2_tiehi
X_09086_ net1316 VGND VPWR _01141_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[6\]
+ clknet_leaf_140_clk_regs sg13g2_dfrbpq_1
X_05318_ net1110 _02038_ _02043_ VPWR VGND sg13g2_nor2_1
X_08106_ net588 VGND VPWR _00187_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[11\]
+ clknet_leaf_125_clk_regs sg13g2_dfrbpq_1
X_08037_ net657 VGND VPWR _00118_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[6\]
+ clknet_leaf_56_clk_regs sg13g2_dfrbpq_1
X_05249_ _01974_ _01975_ net39 VPWR VGND sg13g2_nor2_1
Xhold840 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[22\]
+ VPWR VGND net2667 sg13g2_dlygate4sd3_1
Xhold851 _00732_ VPWR VGND net2678 sg13g2_dlygate4sd3_1
Xhold862 _00707_ VPWR VGND net2689 sg13g2_dlygate4sd3_1
Xhold873 _00239_ VPWR VGND net2700 sg13g2_dlygate4sd3_1
XFILLER_104_944 VPWR VGND sg13g2_decap_8
Xhold895 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[16\]
+ VPWR VGND net2722 sg13g2_dlygate4sd3_1
Xhold884 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[24\]
+ VPWR VGND net2711 sg13g2_dlygate4sd3_1
XFILLER_103_465 VPWR VGND sg13g2_decap_8
XFILLER_67_36 VPWR VGND sg13g2_fill_1
X_08939_ net1463 VGND VPWR net2655 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[5\]
+ clknet_leaf_67_clk_regs sg13g2_dfrbpq_1
Xhold1551 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[11\]
+ VPWR VGND net3378 sg13g2_dlygate4sd3_1
Xhold1540 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[18\]
+ VPWR VGND net3367 sg13g2_dlygate4sd3_1
Xhold1562 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[25\]
+ VPWR VGND net3389 sg13g2_dlygate4sd3_1
XFILLER_29_232 VPWR VGND sg13g2_fill_1
Xhold1573 _02387_ VPWR VGND net3400 sg13g2_dlygate4sd3_1
Xhold1584 i_exotiny._0018_\[0\] VPWR VGND net3411 sg13g2_dlygate4sd3_1
Xhold1595 i_exotiny._1618_\[1\] VPWR VGND net3422 sg13g2_dlygate4sd3_1
XFILLER_26_950 VPWR VGND sg13g2_fill_2
X_08445__236 VPWR VGND net236 sg13g2_tiehi
XFILLER_53_791 VPWR VGND sg13g2_fill_1
Xclkbuf_5_21__f_clk_regs clknet_4_10_0_clk_regs clknet_5_21__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_5_854 VPWR VGND sg13g2_decap_8
XFILLER_80_1028 VPWR VGND sg13g2_fill_1
XFILLER_94_113 VPWR VGND sg13g2_fill_2
XFILLER_94_124 VPWR VGND sg13g2_fill_1
XFILLER_94_179 VPWR VGND sg13g2_fill_1
X_04620_ VPWR _01382_ net1244 VGND sg13g2_inv_1
X_07270_ _02976_ net2614 net1003 _00990_ VPWR VGND sg13g2_mux2_1
XFILLER_32_953 VPWR VGND sg13g2_fill_1
X_06221_ _02542_ net3455 net945 _00375_ VPWR VGND sg13g2_mux2_1
X_06152_ i_exotiny._0028_\[0\] net3127 net953 _00314_ VPWR VGND sg13g2_mux2_1
Xhold103 i_exotiny.i_wb_spi.cnt_hbit_r\[6\] VPWR VGND net1930 sg13g2_dlygate4sd3_1
Xhold114 i_exotiny._1924_\[8\] VPWR VGND net1941 sg13g2_dlygate4sd3_1
Xhold125 _00945_ VPWR VGND net1952 sg13g2_dlygate4sd3_1
X_06083_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[9\]
+ net2148 net955 _00259_ VPWR VGND sg13g2_mux2_1
XFILLER_7_191 VPWR VGND sg13g2_fill_2
X_05103_ _01830_ VPWR _01833_ VGND _01677_ _01815_ sg13g2_o21ai_1
XFILLER_104_229 VPWR VGND sg13g2_decap_8
Xhold136 i_exotiny._1924_\[15\] VPWR VGND net1963 sg13g2_dlygate4sd3_1
Xhold147 i_exotiny._0314_\[27\] VPWR VGND net1974 sg13g2_dlygate4sd3_1
Xhold158 _02254_ VPWR VGND net1985 sg13g2_dlygate4sd3_1
X_05034_ net1220 _01756_ _01759_ _01766_ VPWR VGND sg13g2_nor3_2
Xhold169 i_exotiny._1160_\[5\] VPWR VGND net1996 sg13g2_dlygate4sd3_1
XFILLER_100_402 VPWR VGND sg13g2_decap_8
XFILLER_99_975 VPWR VGND sg13g2_decap_8
XFILLER_98_474 VPWR VGND sg13g2_decap_8
XFILLER_58_305 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_131_clk_regs clknet_5_20__leaf_clk_regs clknet_leaf_131_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_101_969 VPWR VGND sg13g2_decap_8
X_06985_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[27\]
+ net2178 net1019 _00758_ VPWR VGND sg13g2_mux2_1
X_09105__877 VPWR VGND net1297 sg13g2_tiehi
X_08724_ net1684 VGND VPWR net2913 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[19\]
+ clknet_leaf_117_clk_regs sg13g2_dfrbpq_1
XFILLER_100_479 VPWR VGND sg13g2_decap_8
X_05936_ i_exotiny._0020_\[1\] net3029 net969 _00145_ VPWR VGND sg13g2_mux2_1
XFILLER_2_1006 VPWR VGND sg13g2_decap_8
X_05867_ i_exotiny._0018_\[1\] net885 _02421_ _02455_ VPWR VGND sg13g2_mux2_1
X_08655_ net1742 VGND VPWR _00723_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[24\]
+ clknet_leaf_147_clk_regs sg13g2_dfrbpq_1
X_07606_ net3235 _03173_ _03175_ VPWR VGND sg13g2_and2_1
XFILLER_53_27 VPWR VGND sg13g2_fill_2
X_08586_ net740 VGND VPWR _00659_ i_exotiny._0314_\[31\] clknet_leaf_4_clk_regs sg13g2_dfrbpq_1
X_04818_ _01559_ net1265 net1218 VPWR VGND sg13g2_nand2_1
X_05798_ _01472_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_hlt_pc_ccx _01598_ _02415_
+ VPWR VGND sg13g2_a21o_1
X_07537_ VGND VPWR _03128_ _03130_ _01103_ net1196 sg13g2_a21oi_1
X_04749_ net1279 i_exotiny._1623_ _01503_ VPWR VGND sg13g2_and2_1
X_09151__831 VPWR VGND net831 sg13g2_tiehi
X_07468_ _03102_ net1148 _03041_ VPWR VGND sg13g2_nand2_1
X_09207_ net772 VGND VPWR net3051 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[29\]
+ clknet_leaf_79_clk_regs sg13g2_dfrbpq_1
X_06419_ _02595_ net3618 _02599_ _00516_ VPWR VGND sg13g2_a21o_1
X_07399_ _03051_ i_exotiny._1840_\[11\] _02992_ VPWR VGND sg13g2_nand2_1
X_09138_ net844 VGND VPWR net2173 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[26\]
+ clknet_leaf_157_clk_regs sg13g2_dfrbpq_1
X_09069_ net1333 VGND VPWR _01124_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[9\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_2_824 VPWR VGND sg13g2_decap_8
XFILLER_104_741 VPWR VGND sg13g2_decap_8
Xhold681 _00423_ VPWR VGND net2508 sg13g2_dlygate4sd3_1
Xhold670 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[31\]
+ VPWR VGND net2497 sg13g2_dlygate4sd3_1
Xhold692 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[23\]
+ VPWR VGND net2519 sg13g2_dlygate4sd3_1
XFILLER_1_345 VPWR VGND sg13g2_fill_1
XFILLER_103_262 VPWR VGND sg13g2_decap_8
XFILLER_64_308 VPWR VGND sg13g2_fill_1
Xclkbuf_5_5__f_clk_regs clknet_4_2_0_clk_regs clknet_5_5__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_100_980 VPWR VGND sg13g2_decap_8
XFILLER_92_639 VPWR VGND sg13g2_fill_1
Xhold1370 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[17\]
+ VPWR VGND net3197 sg13g2_dlygate4sd3_1
Xhold1392 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[11\]
+ VPWR VGND net3219 sg13g2_dlygate4sd3_1
Xhold1381 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[31\]
+ VPWR VGND net3208 sg13g2_dlygate4sd3_1
XFILLER_45_533 VPWR VGND sg13g2_fill_2
XFILLER_9_412 VPWR VGND sg13g2_fill_1
XFILLER_43_93 VPWR VGND sg13g2_fill_1
X_10677_ _10677_/A net26 VPWR VGND sg13g2_buf_1
XFILLER_99_216 VPWR VGND sg13g2_fill_2
XFILLER_4_32 VPWR VGND sg13g2_fill_2
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_96_956 VPWR VGND sg13g2_decap_8
X_06770_ VGND VPWR _01414_ net1190 _02795_ net1169 sg13g2_a21oi_1
X_09259__243 VPWR VGND net243 sg13g2_tiehi
X_05721_ VGND VPWR i_exotiny._1618_\[2\] net1114 _02362_ _02361_ sg13g2_a21oi_1
X_05652_ net1125 i_exotiny._1924_\[13\] _02310_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_577 VPWR VGND sg13g2_decap_4
X_08440_ net245 VGND VPWR net2015 i_exotiny._0369_\[4\] clknet_leaf_11_clk_regs sg13g2_dfrbpq_2
X_04603_ net3730 _01365_ VPWR VGND sg13g2_inv_4
XFILLER_23_216 VPWR VGND sg13g2_fill_2
XFILLER_24_739 VPWR VGND sg13g2_fill_2
X_08371_ net307 VGND VPWR _00452_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[9\]
+ clknet_leaf_138_clk_regs sg13g2_dfrbpq_1
X_05583_ i_exotiny._0352_ _02257_ net1269 _02258_ VPWR VGND sg13g2_nand3_1
X_07322_ _02987_ VPWR _01031_ VGND _01381_ net1150 sg13g2_o21ai_1
XFILLER_104_1028 VPWR VGND sg13g2_fill_1
X_07253_ net2309 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[16\]
+ net1004 _00976_ VPWR VGND sg13g2_mux2_1
X_06204_ net2863 net3205 net947 _00359_ VPWR VGND sg13g2_mux2_1
X_07184_ net3762 net1233 i_exotiny._0315_\[4\] _02956_ VGND VPWR _02594_ sg13g2_nor4_2
X_06135_ net3011 net2261 net1045 _00304_ VPWR VGND sg13g2_mux2_1
X_06066_ i_exotiny._0025_\[3\] net873 _02510_ _02515_ VPWR VGND sg13g2_mux2_1
X_05017_ _01385_ VPWR _01749_ VGND _01747_ _01748_ sg13g2_o21ai_1
XFILLER_100_210 VPWR VGND sg13g2_decap_4
XFILLER_98_271 VPWR VGND sg13g2_decap_8
XFILLER_48_49 VPWR VGND sg13g2_fill_1
XFILLER_87_978 VPWR VGND sg13g2_decap_8
XFILLER_100_276 VPWR VGND sg13g2_decap_8
X_06968_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[10\]
+ net3216 net1020 _00741_ VPWR VGND sg13g2_mux2_1
X_05919_ net2693 net3120 net975 _00136_ VPWR VGND sg13g2_mux2_1
XFILLER_39_393 VPWR VGND sg13g2_fill_1
X_08707_ net1701 VGND VPWR net2628 i_exotiny._0032_\[2\] clknet_leaf_116_clk_regs
+ sg13g2_dfrbpq_2
X_08638_ net1759 VGND VPWR _00706_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[7\]
+ clknet_leaf_146_clk_regs sg13g2_dfrbpq_1
X_06899_ _02901_ _02719_ _02471_ net1068 net3816 VPWR VGND sg13g2_a22oi_1
XFILLER_81_171 VPWR VGND sg13g2_fill_2
X_08569_ net66 VGND VPWR net3403 i_exotiny._0314_\[14\] clknet_leaf_166_clk_regs sg13g2_dfrbpq_1
XFILLER_11_967 VPWR VGND sg13g2_decap_8
XFILLER_7_905 VPWR VGND sg13g2_decap_8
XFILLER_104_593 VPWR VGND sg13g2_decap_4
Xfanout991 net992 net991 VPWR VGND sg13g2_buf_8
XFILLER_64_116 VPWR VGND sg13g2_fill_2
Xfanout980 _03229_ net980 VPWR VGND sg13g2_buf_8
XFILLER_45_352 VPWR VGND sg13g2_fill_1
XFILLER_72_160 VPWR VGND sg13g2_fill_2
XFILLER_54_92 VPWR VGND sg13g2_fill_2
XFILLER_9_242 VPWR VGND sg13g2_fill_1
XFILLER_14_794 VPWR VGND sg13g2_fill_1
X_08399__683 VPWR VGND net683 sg13g2_tiehi
Xclkload23 clkload23/Y clknet_leaf_28_clk_regs VPWR VGND sg13g2_inv_2
Xclkload34 VPWR clkload34/Y clknet_leaf_130_clk_regs VGND sg13g2_inv_1
Xclkload12 VPWR clkload12/Y clknet_leaf_11_clk_regs VGND sg13g2_inv_1
X_08553__702 VPWR VGND net702 sg13g2_tiehi
XFILLER_5_470 VPWR VGND sg13g2_fill_2
X_07940_ net1175 VGND VPWR net2034 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.genblk7.g_value.r_value[0]
+ clknet_leaf_37_clk_regs sg13g2_dfrbpq_1
X_07871_ net2365 net2690 net978 _01338_ VPWR VGND sg13g2_mux2_1
X_09141__841 VPWR VGND net841 sg13g2_tiehi
X_06822_ net1170 VPWR _02839_ VGND net3644 net1185 sg13g2_o21ai_1
XFILLER_56_617 VPWR VGND sg13g2_decap_8
XFILLER_83_458 VPWR VGND sg13g2_fill_1
X_06753_ VPWR VGND net2106 _02780_ net3821 net3791 _02781_ net1182 sg13g2_a221oi_1
XFILLER_93_1005 VPWR VGND sg13g2_decap_8
XFILLER_92_970 VPWR VGND sg13g2_decap_8
X_05704_ VGND VPWR i_exotiny._1619_\[2\] net1114 _02349_ _02348_ sg13g2_a21oi_1
X_06684_ _02721_ net1219 VPWR VGND net1181 sg13g2_nand2b_2
XFILLER_36_385 VPWR VGND sg13g2_fill_1
X_05635_ net2006 net1065 _02297_ VPWR VGND sg13g2_nor2_1
X_08423_ net262 VGND VPWR net2197 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[22\]
+ clknet_leaf_97_clk_regs sg13g2_dfrbpq_1
X_08354_ net324 VGND VPWR _00435_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[24\]
+ clknet_leaf_95_clk_regs sg13g2_dfrbpq_1
X_05566_ net1266 VPWR _02247_ VGND net3523 net3677 sg13g2_o21ai_1
X_07305_ net881 net2840 _02978_ _02981_ VPWR VGND sg13g2_mux2_1
Xclkload6 VPWR clkload6/Y clknet_5_31__leaf_clk_regs VGND sg13g2_inv_1
X_08285_ net393 VGND VPWR net2476 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[19\]
+ clknet_leaf_100_clk_regs sg13g2_dfrbpq_1
X_05497_ VGND VPWR net3603 net1279 _02193_ _02192_ sg13g2_a21oi_1
X_07236_ VGND VPWR net1139 _02972_ _02973_ net1166 sg13g2_a21oi_1
XFILLER_106_825 VPWR VGND sg13g2_decap_8
X_07167_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[28\]
+ net2711 net1011 _00915_ VPWR VGND sg13g2_mux2_1
X_06118_ net2539 net2317 net1047 _00287_ VPWR VGND sg13g2_mux2_1
X_09271__79 VPWR VGND net79 sg13g2_tiehi
XFILLER_105_368 VPWR VGND sg13g2_decap_8
XFILLER_59_48 VPWR VGND sg13g2_fill_2
X_07098_ net3464 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[30\]
+ net917 _00853_ VPWR VGND sg13g2_mux2_1
Xfanout1219 _01447_ net1219 VPWR VGND sg13g2_buf_8
X_06049_ net2391 net2953 net961 _00234_ VPWR VGND sg13g2_mux2_1
Xfanout1208 net1209 net1208 VPWR VGND sg13g2_buf_8
XFILLER_59_455 VPWR VGND sg13g2_decap_4
XFILLER_47_639 VPWR VGND sg13g2_fill_2
X_08915__1067 VPWR VGND net1487 sg13g2_tiehi
XFILLER_43_889 VPWR VGND sg13g2_fill_1
XFILLER_10_241 VPWR VGND sg13g2_fill_2
XFILLER_40_50 VPWR VGND sg13g2_fill_2
XFILLER_40_83 VPWR VGND sg13g2_fill_1
XFILLER_3_963 VPWR VGND sg13g2_decap_8
XFILLER_104_390 VPWR VGND sg13g2_decap_8
XFILLER_78_753 VPWR VGND sg13g2_fill_2
XFILLER_93_701 VPWR VGND sg13g2_fill_2
XFILLER_92_277 VPWR VGND sg13g2_decap_8
X_07987__128 VPWR VGND net128 sg13g2_tiehi
X_05420_ VPWR _02129_ _02128_ VGND sg13g2_inv_1
X_05351_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set[0]
+ net1832 _02073_ VPWR VGND sg13g2_nor2b_1
XFILLER_14_1028 VPWR VGND sg13g2_fill_1
X_08070_ net624 VGND VPWR _00151_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[7\]
+ clknet_leaf_93_clk_regs sg13g2_dfrbpq_1
X_05282_ _02006_ _02007_ _02005_ _02008_ VPWR VGND sg13g2_nand3_1
X_07021_ net2994 net3175 net920 _00788_ VPWR VGND sg13g2_mux2_1
XFILLER_88_506 VPWR VGND sg13g2_fill_1
XFILLER_103_839 VPWR VGND sg13g2_decap_8
XFILLER_69_720 VPWR VGND sg13g2_decap_8
X_08972_ net1430 VGND VPWR _01030_ i_exotiny._0601_ clknet_leaf_10_clk_regs sg13g2_dfrbpq_1
Xhold18 i_exotiny.i_wb_spi.state_r\[23\] VPWR VGND net1845 sg13g2_dlygate4sd3_1
Xhold29 i_exotiny.i_wb_spi.state_r\[22\] VPWR VGND net1856 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_38_clk_regs clknet_5_10__leaf_clk_regs clknet_leaf_38_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_69_764 VPWR VGND sg13g2_fill_2
X_07923_ net725 VGND VPWR net2005 i_exotiny._1924_\[16\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
Xhold1936 i_exotiny.i_rstctl.cnt\[4\] VPWR VGND net3763 sg13g2_dlygate4sd3_1
Xhold1925 _02403_ VPWR VGND net3752 sg13g2_dlygate4sd3_1
Xhold1914 i_exotiny.gpo\[1\] VPWR VGND net3741 sg13g2_dlygate4sd3_1
X_07854_ i_exotiny._0022_\[1\] net882 _03222_ _03225_ VPWR VGND sg13g2_mux2_1
Xhold1903 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data[0]
+ VPWR VGND net3730 sg13g2_dlygate4sd3_1
Xhold1969 _02401_ VPWR VGND net3796 sg13g2_dlygate4sd3_1
Xhold1958 i_exotiny.i_wdg_top.o_wb_dat\[4\] VPWR VGND net3785 sg13g2_dlygate4sd3_1
X_06805_ VGND VPWR _02822_ _02824_ _02825_ net1130 sg13g2_a21oi_1
Xhold1947 _00925_ VPWR VGND net3774 sg13g2_dlygate4sd3_1
X_07950__706 VPWR VGND net706 sg13g2_tiehi
X_07785_ _03216_ net1138 net1165 _03217_ VPWR VGND sg13g2_a21o_2
X_04997_ _01727_ _01728_ _01729_ VPWR VGND sg13g2_and2_1
X_06736_ VGND VPWR net1101 _02765_ _00666_ _02766_ sg13g2_a21oi_1
XFILLER_25_812 VPWR VGND sg13g2_fill_1
XFILLER_37_683 VPWR VGND sg13g2_decap_8
X_06667_ VGND VPWR net3730 _02690_ _02706_ net1153 sg13g2_a21oi_1
X_08406_ net279 VGND VPWR net3262 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[5\]
+ clknet_leaf_90_clk_regs sg13g2_dfrbpq_1
X_05618_ VGND VPWR net1061 _02284_ _00030_ _02282_ sg13g2_a21oi_1
X_06598_ i_exotiny._0314_\[12\] net1159 _02655_ VPWR VGND sg13g2_nor2_1
X_08337_ net341 VGND VPWR _00418_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[7\]
+ clknet_leaf_98_clk_regs sg13g2_dfrbpq_1
XFILLER_20_561 VPWR VGND sg13g2_fill_2
X_05549_ _01553_ _02220_ _02233_ _02234_ VPWR VGND sg13g2_nor3_1
X_08268_ net410 VGND VPWR _00349_ i_exotiny._0033_\[2\] clknet_leaf_102_clk_regs sg13g2_dfrbpq_2
X_07219_ VGND VPWR _01417_ net1090 _00945_ _02970_ sg13g2_a21oi_1
XFILLER_106_622 VPWR VGND sg13g2_decap_8
X_08199_ net478 VGND VPWR net2757 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[30\]
+ clknet_leaf_68_clk_regs sg13g2_dfrbpq_1
XFILLER_10_42 VPWR VGND sg13g2_fill_2
XFILLER_106_699 VPWR VGND sg13g2_decap_8
XFILLER_105_165 VPWR VGND sg13g2_decap_8
Xfanout1016 _02935_ net1016 VPWR VGND sg13g2_buf_8
Xfanout1038 net1042 net1038 VPWR VGND sg13g2_buf_8
Xfanout1027 _02615_ net1027 VPWR VGND sg13g2_buf_8
Xfanout1005 net1006 net1005 VPWR VGND sg13g2_buf_8
XFILLER_0_966 VPWR VGND sg13g2_decap_8
XFILLER_59_252 VPWR VGND sg13g2_fill_1
Xfanout1049 net1052 net1049 VPWR VGND sg13g2_buf_8
XFILLER_87_594 VPWR VGND sg13g2_fill_2
XFILLER_19_84 VPWR VGND sg13g2_fill_1
XFILLER_47_469 VPWR VGND sg13g2_fill_1
XFILLER_34_119 VPWR VGND sg13g2_fill_1
XFILLER_15_322 VPWR VGND sg13g2_fill_2
XFILLER_15_377 VPWR VGND sg13g2_fill_1
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_11_550 VPWR VGND sg13g2_fill_1
X_09131__851 VPWR VGND net851 sg13g2_tiehi
XFILLER_97_303 VPWR VGND sg13g2_decap_8
XFILLER_3_760 VPWR VGND sg13g2_decap_8
XFILLER_2_281 VPWR VGND sg13g2_fill_2
X_04920_ net1255 _01617_ _01640_ _01652_ VPWR VGND sg13g2_nor3_1
X_04851_ _01588_ i_exotiny.i_wb_spi.cnt_presc_r\[3\] _01572_ VPWR VGND sg13g2_xnor2_1
X_07570_ net1225 _01487_ _03151_ net3700 _01114_ VPWR VGND sg13g2_nor4_1
X_04782_ net1246 net1244 _01532_ VPWR VGND sg13g2_nor2_1
X_06521_ net2824 net2902 net929 _00596_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_156_clk_regs clknet_5_19__leaf_clk_regs clknet_leaf_156_clk_regs VPWR
+ VGND sg13g2_buf_8
X_09240_ net567 VGND VPWR net2705 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[30\]
+ clknet_leaf_135_clk_regs sg13g2_dfrbpq_1
X_06452_ net2955 net2381 net934 _00539_ VPWR VGND sg13g2_mux2_1
X_05403_ _02117_ i_exotiny._2034_\[5\] _02115_ VPWR VGND sg13g2_xnor2_1
X_09171_ net811 VGND VPWR _01226_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[27\]
+ clknet_leaf_173_clk_regs sg13g2_dfrbpq_1
X_06383_ VGND VPWR net3702 net10 _02573_ net1225 sg13g2_a21oi_1
X_05334_ _02058_ _01912_ _02052_ _02057_ VPWR VGND sg13g2_and3_1
X_08122_ net572 VGND VPWR net2631 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[27\]
+ clknet_leaf_123_clk_regs sg13g2_dfrbpq_1
X_08053_ net641 VGND VPWR _00134_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[22\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
X_07004_ net2765 net2872 net922 _00771_ VPWR VGND sg13g2_mux2_1
X_05265_ _01991_ _01777_ i_exotiny._0013_\[0\] _01770_ i_exotiny._0025_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_05196_ _01924_ i_exotiny._0035_\[1\] _01778_ VPWR VGND sg13g2_nand2_1
Xoutput19 net19 uio_oe[1] VPWR VGND sg13g2_buf_1
XFILLER_103_614 VPWR VGND sg13g2_fill_1
XFILLER_89_837 VPWR VGND sg13g2_fill_1
X_08955_ net1447 VGND VPWR net2104 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[21\]
+ clknet_leaf_54_clk_regs sg13g2_dfrbpq_1
XFILLER_102_168 VPWR VGND sg13g2_decap_8
XFILLER_97_870 VPWR VGND sg13g2_decap_8
X_07906_ i_exotiny._0000_ VGND VPWR net1105 i_exotiny.i_wdg_top.fsm_inst.sw_trg_s1wto
+ clknet_leaf_40_clk_regs sg13g2_dfrbpq_2
XFILLER_69_572 VPWR VGND sg13g2_fill_2
Xhold1711 _01076_ VPWR VGND net3538 sg13g2_dlygate4sd3_1
Xhold1700 _01048_ VPWR VGND net3527 sg13g2_dlygate4sd3_1
Xhold1744 i_exotiny.i_rstctl.sys_res_n VPWR VGND net3571 sg13g2_dlygate4sd3_1
Xhold1733 _00212_ VPWR VGND net3560 sg13g2_dlygate4sd3_1
X_08886_ net1516 VGND VPWR _00944_ i_exotiny.i_wb_spi.dat_rx_r\[16\] clknet_leaf_59_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_5_1015 VPWR VGND sg13g2_decap_8
Xhold1722 i_exotiny._0315_\[18\] VPWR VGND net3549 sg13g2_dlygate4sd3_1
Xhold1766 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[5\]
+ VPWR VGND net3593 sg13g2_dlygate4sd3_1
Xhold1755 i_exotiny.i_wb_spi.dat_rx_r\[30\] VPWR VGND net3582 sg13g2_dlygate4sd3_1
Xhold1777 _00629_ VPWR VGND net3604 sg13g2_dlygate4sd3_1
X_07837_ net3254 net3333 net986 _01310_ VPWR VGND sg13g2_mux2_1
X_07768_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[24\]
+ net2837 net992 _01253_ VPWR VGND sg13g2_mux2_1
Xhold1788 _00686_ VPWR VGND net3615 sg13g2_dlygate4sd3_1
Xhold1799 i_exotiny._0315_\[11\] VPWR VGND net3626 sg13g2_dlygate4sd3_1
X_06719_ VGND VPWR net1102 _02751_ _00663_ _02752_ sg13g2_a21oi_1
XFILLER_53_973 VPWR VGND sg13g2_fill_1
X_07699_ net3009 net873 _03193_ _03198_ VPWR VGND sg13g2_mux2_1
Xclkbuf_5_20__f_clk_regs clknet_4_10_0_clk_regs clknet_5_20__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_12_347 VPWR VGND sg13g2_fill_1
XFILLER_4_546 VPWR VGND sg13g2_decap_8
XFILLER_106_496 VPWR VGND sg13g2_decap_8
XFILLER_97_67 VPWR VGND sg13g2_fill_1
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_102_680 VPWR VGND sg13g2_fill_2
XFILLER_75_531 VPWR VGND sg13g2_fill_2
XFILLER_62_203 VPWR VGND sg13g2_fill_2
XFILLER_62_236 VPWR VGND sg13g2_fill_2
X_08652__1325 VPWR VGND net1745 sg13g2_tiehi
XFILLER_16_675 VPWR VGND sg13g2_fill_2
X_08798__1190 VPWR VGND net1610 sg13g2_tiehi
XFILLER_11_1009 VPWR VGND sg13g2_decap_8
Xhold307 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[4\]
+ VPWR VGND net2134 sg13g2_dlygate4sd3_1
X_08177__500 VPWR VGND net500 sg13g2_tiehi
Xhold329 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[30\]
+ VPWR VGND net2156 sg13g2_dlygate4sd3_1
Xhold318 _00836_ VPWR VGND net2145 sg13g2_dlygate4sd3_1
X_05050_ i_exotiny._0079_\[2\] i_exotiny._0079_\[3\] net1235 _01782_ VGND VPWR _01753_
+ sg13g2_nor4_2
X_08874__1108 VPWR VGND net1528 sg13g2_tiehi
X_08910__1072 VPWR VGND net1492 sg13g2_tiehi
XFILLER_97_155 VPWR VGND sg13g2_fill_1
X_08740_ net1668 VGND VPWR _00798_ i_exotiny._0017_\[3\] clknet_leaf_82_clk_regs sg13g2_dfrbpq_2
X_05952_ net2170 net3424 net970 _00161_ VPWR VGND sg13g2_mux2_1
Xhold1018 _00262_ VPWR VGND net2845 sg13g2_dlygate4sd3_1
Xhold1029 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[9\]
+ VPWR VGND net2856 sg13g2_dlygate4sd3_1
Xhold1007 _01274_ VPWR VGND net2834 sg13g2_dlygate4sd3_1
X_08671_ net1203 VGND VPWR i_exotiny._2043_\[8\] i_exotiny._2034_\[8\] net1229 sg13g2_dfrbpq_2
X_05883_ _02468_ VPWR _02469_ VGND _01498_ _01834_ sg13g2_o21ai_1
XFILLER_38_233 VPWR VGND sg13g2_fill_1
X_04903_ _01635_ i_exotiny._0013_\[3\] _01634_ VPWR VGND sg13g2_nand2_1
X_07622_ VGND VPWR net1228 _03183_ _03185_ net1205 sg13g2_a21oi_1
X_04834_ i_exotiny.i_wb_spi.cnt_presc_r\[4\] _01573_ _01574_ VPWR VGND sg13g2_nor2b_1
X_07553_ _03134_ VPWR _03141_ VGND net3763 _03139_ sg13g2_o21ai_1
X_04765_ net1219 net1181 _01516_ VPWR VGND sg13g2_nor2_1
X_06504_ _02617_ net2532 net1025 _00583_ VPWR VGND sg13g2_mux2_1
X_07484_ _03109_ net1233 net906 VPWR VGND sg13g2_nand2_1
X_04696_ net1270 _01453_ _01454_ VPWR VGND sg13g2_and2_1
X_06435_ net2905 i_exotiny._0039_\[0\] net938 _00522_ VPWR VGND sg13g2_mux2_1
X_09223_ net756 VGND VPWR _01278_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[13\]
+ clknet_leaf_129_clk_regs sg13g2_dfrbpq_1
X_09154_ net828 VGND VPWR net3272 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[10\]
+ clknet_leaf_148_clk_regs sg13g2_dfrbpq_1
X_06366_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[25\]
+ net2473 net1031 _00496_ VPWR VGND sg13g2_mux2_1
X_08105_ net589 VGND VPWR net2378 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[10\]
+ clknet_leaf_122_clk_regs sg13g2_dfrbpq_1
X_06297_ _02554_ net2383 net941 _00439_ VPWR VGND sg13g2_mux2_1
X_09085_ net1317 VGND VPWR _01140_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[5\]
+ clknet_leaf_142_clk_regs sg13g2_dfrbpq_1
X_05317_ _01608_ _02038_ _02042_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_53_clk_regs clknet_5_15__leaf_clk_regs clknet_leaf_53_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08036_ net658 VGND VPWR _00117_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[5\]
+ clknet_leaf_55_clk_regs sg13g2_dfrbpq_1
X_08297__381 VPWR VGND net381 sg13g2_tiehi
Xhold830 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[27\]
+ VPWR VGND net2657 sg13g2_dlygate4sd3_1
X_05248_ VPWR VGND _01944_ net1109 _01920_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[1\]
+ _01975_ net1107 sg13g2_a221oi_1
XFILLER_104_923 VPWR VGND sg13g2_decap_8
Xhold841 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[27\]
+ VPWR VGND net2668 sg13g2_dlygate4sd3_1
Xhold863 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[13\]
+ VPWR VGND net2690 sg13g2_dlygate4sd3_1
Xhold852 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[19\]
+ VPWR VGND net2679 sg13g2_dlygate4sd3_1
Xhold896 _00743_ VPWR VGND net2723 sg13g2_dlygate4sd3_1
Xhold874 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[20\]
+ VPWR VGND net2701 sg13g2_dlygate4sd3_1
Xhold885 _00915_ VPWR VGND net2712 sg13g2_dlygate4sd3_1
X_05179_ _01831_ _01902_ _01903_ _01907_ VPWR VGND sg13g2_or3_1
XFILLER_103_444 VPWR VGND sg13g2_decap_8
Xclkbuf_5_4__f_clk_regs clknet_4_2_0_clk_regs clknet_5_4__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08730__1258 VPWR VGND net1678 sg13g2_tiehi
X_08938_ net1464 VGND VPWR _00996_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[4\]
+ clknet_leaf_74_clk_regs sg13g2_dfrbpq_1
Xhold1530 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[23\]
+ VPWR VGND net3357 sg13g2_dlygate4sd3_1
Xhold1552 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[9\]
+ VPWR VGND net3379 sg13g2_dlygate4sd3_1
X_08869_ net1534 VGND VPWR net3746 i_exotiny.gpo\[2\] clknet_leaf_29_clk_regs sg13g2_dfrbpq_1
XFILLER_18_918 VPWR VGND sg13g2_fill_1
Xhold1541 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[5\]
+ VPWR VGND net3368 sg13g2_dlygate4sd3_1
Xhold1574 _00064_ VPWR VGND net3401 sg13g2_dlygate4sd3_1
Xhold1585 i_exotiny._0038_\[3\] VPWR VGND net3412 sg13g2_dlygate4sd3_1
X_09121__861 VPWR VGND net861 sg13g2_tiehi
Xhold1563 i_exotiny._0314_\[3\] VPWR VGND net3390 sg13g2_dlygate4sd3_1
XFILLER_29_255 VPWR VGND sg13g2_fill_1
Xhold1596 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[12\]
+ VPWR VGND net3423 sg13g2_dlygate4sd3_1
XFILLER_41_910 VPWR VGND sg13g2_decap_4
XFILLER_41_965 VPWR VGND sg13g2_fill_1
XFILLER_5_833 VPWR VGND sg13g2_decap_8
XFILLER_5_811 VPWR VGND sg13g2_decap_4
XFILLER_5_800 VPWR VGND sg13g2_fill_2
XFILLER_99_409 VPWR VGND sg13g2_decap_8
XFILLER_106_293 VPWR VGND sg13g2_decap_8
X_08706__1282 VPWR VGND net1702 sg13g2_tiehi
X_09237__701 VPWR VGND net701 sg13g2_tiehi
XFILLER_90_353 VPWR VGND sg13g2_fill_1
X_08601__1375 VPWR VGND net1795 sg13g2_tiehi
X_06220_ i_exotiny._0033_\[0\] net888 _02540_ _02542_ VPWR VGND sg13g2_mux2_1
X_08928__1054 VPWR VGND net1474 sg13g2_tiehi
X_06151_ net1158 VPWR _02534_ VGND _02423_ _02533_ sg13g2_o21ai_1
Xhold104 _02380_ VPWR VGND net1931 sg13g2_dlygate4sd3_1
Xhold126 i_exotiny._1924_\[13\] VPWR VGND net1953 sg13g2_dlygate4sd3_1
Xhold115 _00033_ VPWR VGND net1942 sg13g2_dlygate4sd3_1
X_06082_ net3349 net3423 net955 _00258_ VPWR VGND sg13g2_mux2_1
XFILLER_7_170 VPWR VGND sg13g2_fill_1
X_08537__143 VPWR VGND net143 sg13g2_tiehi
X_05102_ _01677_ _01815_ _01830_ _01832_ VPWR VGND sg13g2_or3_1
XFILLER_104_208 VPWR VGND sg13g2_decap_8
Xhold137 _00040_ VPWR VGND net1964 sg13g2_dlygate4sd3_1
Xhold148 _00651_ VPWR VGND net1975 sg13g2_dlygate4sd3_1
Xhold159 i_exotiny._1489_\[2\] VPWR VGND net1986 sg13g2_dlygate4sd3_1
X_05033_ net1220 _01753_ _01757_ _01765_ VPWR VGND sg13g2_nor3_2
XFILLER_99_954 VPWR VGND sg13g2_decap_8
XFILLER_98_453 VPWR VGND sg13g2_decap_8
XFILLER_101_948 VPWR VGND sg13g2_decap_8
X_06984_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[26\]
+ net2160 net1020 _00757_ VPWR VGND sg13g2_mux2_1
XFILLER_100_458 VPWR VGND sg13g2_decap_8
X_05935_ i_exotiny._0020_\[0\] net2675 net968 _00144_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_171_clk_regs clknet_5_5__leaf_clk_regs clknet_leaf_171_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08723_ net1685 VGND VPWR _00781_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[18\]
+ clknet_leaf_121_clk_regs sg13g2_dfrbpq_1
XFILLER_73_309 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_100_clk_regs clknet_5_29__leaf_clk_regs clknet_leaf_100_clk_regs VPWR
+ VGND sg13g2_buf_8
X_05866_ _01470_ _02453_ _02454_ VPWR VGND sg13g2_nor2_2
X_08654_ net1743 VGND VPWR _00722_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[23\]
+ clknet_leaf_146_clk_regs sg13g2_dfrbpq_1
X_07605_ net3235 _03173_ _03174_ VPWR VGND sg13g2_nor2_1
X_04817_ net19 _01557_ _01558_ VPWR VGND sg13g2_nand2_2
X_08585_ net1812 VGND VPWR net3731 i_exotiny._0314_\[30\] clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
XFILLER_26_269 VPWR VGND sg13g2_fill_2
X_05797_ VGND VPWR _01598_ _02414_ _01472_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_hlt_pc_ccx
+ sg13g2_a21oi_2
XFILLER_42_707 VPWR VGND sg13g2_fill_1
XFILLER_42_718 VPWR VGND sg13g2_fill_1
X_04748_ i_exotiny._1265_ _01465_ net1268 _01502_ VPWR VGND sg13g2_nand3_1
X_07536_ _03126_ _03129_ _01442_ _03130_ VPWR VGND sg13g2_nand3_1
X_09206_ net773 VGND VPWR net3008 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[28\]
+ clknet_leaf_78_clk_regs sg13g2_dfrbpq_1
X_04679_ _01439_ net3827 _01440_ VPWR VGND sg13g2_xor2_1
X_07467_ net1207 _02989_ net3415 _03101_ VPWR VGND sg13g2_nand3_1
X_06418_ net1282 VPWR _02599_ VGND _01366_ _02595_ sg13g2_o21ai_1
X_07398_ _03050_ _02992_ _02998_ VPWR VGND sg13g2_nand2_1
X_06349_ net2929 net2138 net1029 _00479_ VPWR VGND sg13g2_mux2_1
X_09137_ net845 VGND VPWR net2728 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[25\]
+ clknet_leaf_154_clk_regs sg13g2_dfrbpq_1
X_09068_ net1334 VGND VPWR _01123_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[8\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_1
X_08019_ net675 VGND VPWR _00100_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[20\]
+ clknet_leaf_62_clk_regs sg13g2_dfrbpq_1
XFILLER_2_803 VPWR VGND sg13g2_decap_8
XFILLER_104_720 VPWR VGND sg13g2_decap_8
Xhold660 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[14\]
+ VPWR VGND net2487 sg13g2_dlygate4sd3_1
Xhold671 _01292_ VPWR VGND net2498 sg13g2_dlygate4sd3_1
XFILLER_103_241 VPWR VGND sg13g2_decap_8
Xhold682 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[30\]
+ VPWR VGND net2509 sg13g2_dlygate4sd3_1
Xhold693 _01256_ VPWR VGND net2520 sg13g2_dlygate4sd3_1
XFILLER_89_464 VPWR VGND sg13g2_fill_2
XFILLER_89_453 VPWR VGND sg13g2_fill_1
XFILLER_89_442 VPWR VGND sg13g2_fill_1
XFILLER_104_797 VPWR VGND sg13g2_decap_8
Xhold1360 i_exotiny._0029_\[1\] VPWR VGND net3187 sg13g2_dlygate4sd3_1
X_08564__76 VPWR VGND net76 sg13g2_tiehi
Xhold1382 _00378_ VPWR VGND net3209 sg13g2_dlygate4sd3_1
Xhold1371 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[15\]
+ VPWR VGND net3198 sg13g2_dlygate4sd3_1
Xhold1393 i_exotiny._0315_\[25\] VPWR VGND net3220 sg13g2_dlygate4sd3_1
XFILLER_26_792 VPWR VGND sg13g2_fill_1
XFILLER_14_943 VPWR VGND sg13g2_fill_2
XFILLER_41_784 VPWR VGND sg13g2_fill_1
X_10676_ i_exotiny.i_wb_spi.spi_sdo_o net25 VPWR VGND sg13g2_buf_1
XFILLER_99_206 VPWR VGND sg13g2_fill_1
X_08174__503 VPWR VGND net503 sg13g2_tiehi
X_08619__1357 VPWR VGND net1777 sg13g2_tiehi
XFILLER_96_935 VPWR VGND sg13g2_decap_8
XFILLER_1_880 VPWR VGND sg13g2_decap_8
XFILLER_95_434 VPWR VGND sg13g2_decap_4
X_09204__777 VPWR VGND net777 sg13g2_tiehi
X_05720_ net1114 i_exotiny._1924_\[30\] _02361_ VPWR VGND sg13g2_nor2b_1
X_05651_ net1939 net1066 _02309_ VPWR VGND sg13g2_nor2_1
XFILLER_63_342 VPWR VGND sg13g2_fill_1
X_08287__391 VPWR VGND net391 sg13g2_tiehi
X_04602_ VPWR _01364_ i_exotiny.gpo\[2\] VGND sg13g2_inv_1
X_08370_ net308 VGND VPWR _00451_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[8\]
+ clknet_leaf_137_clk_regs sg13g2_dfrbpq_1
X_05582_ _01465_ net1201 _02257_ VPWR VGND _01461_ sg13g2_nand3b_1
X_07321_ _02987_ net3643 net1151 VPWR VGND sg13g2_nand2_1
XFILLER_104_1007 VPWR VGND sg13g2_decap_8
X_07252_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[19\]
+ net3352 net1006 _00975_ VPWR VGND sg13g2_mux2_1
X_07183_ _00924_ _02954_ net2107 _02953_ _01367_ VPWR VGND sg13g2_a22oi_1
X_06203_ net3479 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[11\]
+ net949 _00358_ VPWR VGND sg13g2_mux2_1
X_09283__55 VPWR VGND net55 sg13g2_tiehi
X_06134_ net2389 net3171 net1047 _00303_ VPWR VGND sg13g2_mux2_1
X_09111__871 VPWR VGND net871 sg13g2_tiehi
X_06065_ _02514_ net2271 net962 _00247_ VPWR VGND sg13g2_mux2_1
XFILLER_98_250 VPWR VGND sg13g2_decap_8
X_08294__384 VPWR VGND net384 sg13g2_tiehi
X_05016_ _01746_ _01729_ _01701_ _01748_ VPWR VGND sg13g2_a21o_1
XFILLER_100_255 VPWR VGND sg13g2_decap_8
XFILLER_55_810 VPWR VGND sg13g2_fill_1
X_06967_ net2944 net2988 net1018 _00740_ VPWR VGND sg13g2_mux2_1
X_05918_ net2433 net2668 net973 _00135_ VPWR VGND sg13g2_mux2_1
XFILLER_73_139 VPWR VGND sg13g2_fill_2
XFILLER_66_180 VPWR VGND sg13g2_fill_1
X_06898_ VPWR _00694_ _02900_ VGND sg13g2_inv_1
X_08706_ net1702 VGND VPWR _00764_ i_exotiny._0032_\[1\] clknet_leaf_116_clk_regs
+ sg13g2_dfrbpq_2
X_08637_ net1760 VGND VPWR _00705_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[6\]
+ clknet_leaf_150_clk_regs sg13g2_dfrbpq_1
X_05849_ _02438_ _02437_ _01470_ VPWR VGND sg13g2_nand2b_1
X_08568_ net68 VGND VPWR net2865 i_exotiny._0314_\[13\] clknet_leaf_180_clk_regs sg13g2_dfrbpq_1
XFILLER_70_1028 VPWR VGND sg13g2_fill_1
X_08499_ net181 VGND VPWR net2941 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[19\]
+ clknet_leaf_107_clk_regs sg13g2_dfrbpq_1
X_07519_ _01945_ _01499_ net901 _03117_ VPWR VGND sg13g2_a21o_1
XFILLER_50_592 VPWR VGND sg13g2_fill_2
XFILLER_11_946 VPWR VGND sg13g2_decap_8
XFILLER_22_294 VPWR VGND sg13g2_fill_1
XFILLER_8_2 VPWR VGND sg13g2_fill_1
Xhold490 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[5\]
+ VPWR VGND net2317 sg13g2_dlygate4sd3_1
XFILLER_1_154 VPWR VGND sg13g2_fill_1
XFILLER_93_905 VPWR VGND sg13g2_fill_1
Xfanout970 net971 net970 VPWR VGND sg13g2_buf_2
Xfanout992 _03211_ net992 VPWR VGND sg13g2_buf_8
XFILLER_93_949 VPWR VGND sg13g2_decap_8
Xfanout981 net982 net981 VPWR VGND sg13g2_buf_8
XFILLER_46_810 VPWR VGND sg13g2_fill_1
XFILLER_86_990 VPWR VGND sg13g2_decap_8
XFILLER_38_94 VPWR VGND sg13g2_fill_2
Xhold1190 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[28\]
+ VPWR VGND net3017 sg13g2_dlygate4sd3_1
X_08527__153 VPWR VGND net153 sg13g2_tiehi
XFILLER_60_334 VPWR VGND sg13g2_fill_2
XFILLER_20_209 VPWR VGND sg13g2_fill_1
Xclkload24 clkload24/Y clknet_leaf_36_clk_regs VPWR VGND sg13g2_inv_2
Xclkload35 clkload35/Y clknet_leaf_136_clk_regs VPWR VGND sg13g2_inv_2
X_09265__99 VPWR VGND net99 sg13g2_tiehi
Xclkload13 clkload13/Y clknet_leaf_12_clk_regs VPWR VGND sg13g2_inv_2
XFILLER_6_983 VPWR VGND sg13g2_decap_8
X_08534__146 VPWR VGND net146 sg13g2_tiehi
XFILLER_69_935 VPWR VGND sg13g2_fill_2
XFILLER_69_924 VPWR VGND sg13g2_fill_1
XFILLER_69_968 VPWR VGND sg13g2_fill_2
X_07870_ net2684 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[12\]
+ net979 _01337_ VPWR VGND sg13g2_mux2_1
X_06821_ i_exotiny._0369_\[20\] net1188 _02838_ VPWR VGND sg13g2_nor2_1
XFILLER_95_286 VPWR VGND sg13g2_decap_8
X_06752_ VGND VPWR _01406_ _01451_ _02780_ _02779_ sg13g2_a21oi_1
X_05703_ net1115 i_exotiny._1924_\[26\] _02348_ VPWR VGND sg13g2_nor2b_1
XFILLER_52_802 VPWR VGND sg13g2_fill_2
XFILLER_37_865 VPWR VGND sg13g2_fill_2
XFILLER_93_1028 VPWR VGND sg13g2_fill_1
X_08422_ net263 VGND VPWR net2474 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[21\]
+ clknet_leaf_90_clk_regs sg13g2_dfrbpq_1
X_06683_ _02720_ net1137 net1102 VPWR VGND sg13g2_nand2_1
XFILLER_52_835 VPWR VGND sg13g2_fill_1
X_05634_ VGND VPWR net1066 _02296_ _00034_ _02294_ sg13g2_a21oi_1
X_08541__139 VPWR VGND net139 sg13g2_tiehi
X_08353_ net325 VGND VPWR _00434_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[23\]
+ clknet_leaf_97_clk_regs sg13g2_dfrbpq_1
XFILLER_51_378 VPWR VGND sg13g2_fill_1
X_05565_ VGND VPWR net1202 _02244_ _02246_ _02245_ sg13g2_a21oi_1
X_07304_ net3232 _02980_ net909 _01020_ VPWR VGND sg13g2_mux2_1
X_08284_ net394 VGND VPWR net2567 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[18\]
+ clknet_leaf_103_clk_regs sg13g2_dfrbpq_1
X_07235_ _02518_ _02564_ _02972_ VPWR VGND sg13g2_nor2_2
Xclkload7 clknet_leaf_186_clk_regs clkload7/X VPWR VGND sg13g2_buf_8
X_05496_ net1279 _01393_ _02192_ VPWR VGND sg13g2_nor2_1
XFILLER_106_804 VPWR VGND sg13g2_decap_8
X_07166_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[27\]
+ net2442 net1009 _00914_ VPWR VGND sg13g2_mux2_1
X_06117_ net2762 net3111 net1043 _00286_ VPWR VGND sg13g2_mux2_1
X_07097_ net2512 net2936 net913 _00852_ VPWR VGND sg13g2_mux2_1
XFILLER_105_347 VPWR VGND sg13g2_decap_8
X_06048_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[20\]
+ net2220 net965 _00233_ VPWR VGND sg13g2_mux2_1
Xfanout1209 net1210 net1209 VPWR VGND sg13g2_buf_8
XFILLER_101_520 VPWR VGND sg13g2_decap_4
X_07999_ net696 VGND VPWR net2485 i_exotiny._0018_\[0\] clknet_leaf_67_clk_regs sg13g2_dfrbpq_2
XFILLER_27_320 VPWR VGND sg13g2_fill_1
XFILLER_54_172 VPWR VGND sg13g2_fill_2
XFILLER_70_632 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_8_clk_regs clknet_5_2__leaf_clk_regs clknet_leaf_8_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_6_268 VPWR VGND sg13g2_fill_2
XFILLER_3_942 VPWR VGND sg13g2_decap_8
XFILLER_105_881 VPWR VGND sg13g2_decap_8
X_08171__506 VPWR VGND net506 sg13g2_tiehi
XFILLER_1_56 VPWR VGND sg13g2_fill_2
XFILLER_92_256 VPWR VGND sg13g2_fill_2
X_08743__1245 VPWR VGND net1665 sg13g2_tiehi
XFILLER_65_70 VPWR VGND sg13g2_fill_1
X_09101__881 VPWR VGND net1301 sg13g2_tiehi
XFILLER_34_835 VPWR VGND sg13g2_fill_1
X_05350_ net1263 net3780 _02072_ VPWR VGND sg13g2_nor2_1
X_08284__394 VPWR VGND net394 sg13g2_tiehi
XFILLER_33_389 VPWR VGND sg13g2_fill_1
X_05281_ _02007_ _01778_ i_exotiny._0035_\[0\] _01773_ i_exotiny._0019_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_07020_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[24\]
+ net2083 net922 _00787_ VPWR VGND sg13g2_mux2_1
X_08965__1017 VPWR VGND net1437 sg13g2_tiehi
XFILLER_6_780 VPWR VGND sg13g2_decap_4
XFILLER_103_818 VPWR VGND sg13g2_decap_8
X_08971_ net1431 VGND VPWR _01029_ i_exotiny._0542_ clknet_leaf_10_clk_regs sg13g2_dfrbpq_1
Xhold19 i_exotiny.i_wb_spi.state_r\[8\] VPWR VGND net1846 sg13g2_dlygate4sd3_1
X_07922_ net726 VGND VPWR net1964 i_exotiny._1924_\[15\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
Xhold1926 _00072_ VPWR VGND net3753 sg13g2_dlygate4sd3_1
X_08291__387 VPWR VGND net387 sg13g2_tiehi
XFILLER_57_905 VPWR VGND sg13g2_fill_2
Xhold1915 _02958_ VPWR VGND net3742 sg13g2_dlygate4sd3_1
Xhold1904 _00658_ VPWR VGND net3731 sg13g2_dlygate4sd3_1
X_07853_ _03224_ net2471 net985 _01325_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_78_clk_regs clknet_5_26__leaf_clk_regs clknet_leaf_78_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold1959 _00070_ VPWR VGND net3786 sg13g2_dlygate4sd3_1
XFILLER_68_286 VPWR VGND sg13g2_fill_1
X_06804_ _02823_ VPWR _02824_ VGND net3675 net1191 sg13g2_o21ai_1
XFILLER_56_437 VPWR VGND sg13g2_decap_8
Xhold1948 i_exotiny.i_wb_qspi_mem.crm_r VPWR VGND net3775 sg13g2_dlygate4sd3_1
Xhold1937 i_exotiny._0369_\[28\] VPWR VGND net3764 sg13g2_dlygate4sd3_1
X_07784_ _02485_ _02518_ _03216_ VPWR VGND sg13g2_nor2_2
XFILLER_37_651 VPWR VGND sg13g2_decap_4
X_04996_ _01728_ _01712_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data[0]
+ VPWR VGND sg13g2_nand2b_1
X_06735_ net3730 net1101 _02766_ VPWR VGND sg13g2_nor2_1
XFILLER_52_643 VPWR VGND sg13g2_decap_8
X_06666_ _02705_ _02703_ _02704_ VPWR VGND sg13g2_nand2b_1
X_08405_ net280 VGND VPWR _00479_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[4\]
+ clknet_leaf_94_clk_regs sg13g2_dfrbpq_1
X_05617_ VGND VPWR i_exotiny._1612_\[0\] net1119 _02284_ _02283_ sg13g2_a21oi_1
XFILLER_51_142 VPWR VGND sg13g2_fill_1
XFILLER_51_131 VPWR VGND sg13g2_fill_2
XFILLER_24_367 VPWR VGND sg13g2_fill_2
X_08336_ net342 VGND VPWR _00417_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[6\]
+ clknet_leaf_107_clk_regs sg13g2_dfrbpq_1
X_06597_ net1198 _02653_ _02654_ _00639_ VPWR VGND sg13g2_nor3_1
X_05548_ _02221_ _02232_ _02233_ VPWR VGND sg13g2_nor2_1
X_08614__1362 VPWR VGND net1782 sg13g2_tiehi
X_08267_ net411 VGND VPWR net2231 i_exotiny._0033_\[1\] clknet_leaf_103_clk_regs sg13g2_dfrbpq_2
X_05479_ _02180_ _02178_ _02179_ VPWR VGND sg13g2_nand2_1
XFILLER_106_601 VPWR VGND sg13g2_decap_8
X_07218_ net1951 net1090 _02970_ VPWR VGND sg13g2_nor2_1
X_08198_ net479 VGND VPWR _00279_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[29\]
+ clknet_leaf_112_clk_regs sg13g2_dfrbpq_1
X_07149_ net2787 net3281 net1011 _00897_ VPWR VGND sg13g2_mux2_1
XFILLER_105_144 VPWR VGND sg13g2_decap_8
X_08517__163 VPWR VGND net163 sg13g2_tiehi
XFILLER_106_678 VPWR VGND sg13g2_decap_8
X_08821__1167 VPWR VGND net1587 sg13g2_tiehi
Xfanout1017 _02935_ net1017 VPWR VGND sg13g2_buf_8
Xfanout1028 net1029 net1028 VPWR VGND sg13g2_buf_8
Xfanout1006 net1007 net1006 VPWR VGND sg13g2_buf_8
XFILLER_0_945 VPWR VGND sg13g2_decap_8
Xfanout1039 net1042 net1039 VPWR VGND sg13g2_buf_8
XFILLER_102_895 VPWR VGND sg13g2_decap_8
XFILLER_75_724 VPWR VGND sg13g2_fill_2
XFILLER_101_394 VPWR VGND sg13g2_decap_8
XFILLER_35_51 VPWR VGND sg13g2_decap_4
XFILLER_71_974 VPWR VGND sg13g2_fill_1
X_08524__156 VPWR VGND net156 sg13g2_tiehi
X_08099__595 VPWR VGND net595 sg13g2_tiehi
XFILLER_97_359 VPWR VGND sg13g2_decap_8
X_08531__149 VPWR VGND net149 sg13g2_tiehi
X_04850_ net1111 _01583_ _01587_ i_exotiny._1902_\[2\] VPWR VGND sg13g2_nor3_1
X_04781_ _01529_ _01530_ _01531_ VPWR VGND sg13g2_nor2b_1
X_06520_ net2541 net3132 net932 _00595_ VPWR VGND sg13g2_mux2_1
X_06451_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[20\]
+ net2737 net938 _00538_ VPWR VGND sg13g2_mux2_1
XFILLER_33_142 VPWR VGND sg13g2_fill_2
XFILLER_34_687 VPWR VGND sg13g2_fill_2
X_05402_ net1113 _02115_ _02116_ i_exotiny._2043_\[4\] VPWR VGND sg13g2_nor3_1
XFILLER_33_175 VPWR VGND sg13g2_fill_1
X_09170_ net812 VGND VPWR net2518 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[26\]
+ clknet_leaf_172_clk_regs sg13g2_dfrbpq_1
X_06382_ _02572_ _01524_ _02571_ VPWR VGND sg13g2_nand2_1
X_08121_ net573 VGND VPWR net2157 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[26\]
+ clknet_leaf_122_clk_regs sg13g2_dfrbpq_1
X_05333_ _01818_ _02056_ _02057_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_125_clk_regs clknet_5_23__leaf_clk_regs clknet_leaf_125_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08052_ net642 VGND VPWR net2165 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[21\]
+ clknet_leaf_55_clk_regs sg13g2_dfrbpq_1
X_05264_ _01990_ i_exotiny._0023_\[0\] _01783_ VPWR VGND sg13g2_nand2_1
X_07003_ net2093 net2972 net918 _00770_ VPWR VGND sg13g2_mux2_1
X_05195_ _01923_ _01781_ i_exotiny._0028_\[1\] _01766_ i_exotiny._0030_\[1\] VPWR
+ VGND sg13g2_a22oi_1
X_08954_ net1448 VGND VPWR _01012_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[20\]
+ clknet_leaf_75_clk_regs sg13g2_dfrbpq_1
Xclkbuf_5_3__f_clk_regs clknet_4_1_0_clk_regs clknet_5_3__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold1701 i_exotiny.i_wdg_top.o_wb_dat\[3\] VPWR VGND net3528 sg13g2_dlygate4sd3_1
X_07905_ net1176 VGND VPWR net3568 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.genblk7.g_value.r_value[0]
+ clknet_leaf_38_clk_regs sg13g2_dfrbpq_2
Xhold1712 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[7\]
+ VPWR VGND net3539 sg13g2_dlygate4sd3_1
X_08885_ net1517 VGND VPWR _00943_ i_exotiny.i_wb_spi.dat_rx_r\[15\] clknet_leaf_62_clk_regs
+ sg13g2_dfrbpq_1
Xhold1734 i_exotiny._2025_\[5\] VPWR VGND net3561 sg13g2_dlygate4sd3_1
Xhold1723 _01088_ VPWR VGND net3550 sg13g2_dlygate4sd3_1
XFILLER_96_392 VPWR VGND sg13g2_decap_8
XFILLER_84_532 VPWR VGND sg13g2_fill_1
Xhold1745 i_exotiny._1616_\[1\] VPWR VGND net3572 sg13g2_dlygate4sd3_1
Xhold1756 _00958_ VPWR VGND net3583 sg13g2_dlygate4sd3_1
XFILLER_56_223 VPWR VGND sg13g2_fill_1
Xhold1778 i_exotiny._0314_\[7\] VPWR VGND net3605 sg13g2_dlygate4sd3_1
X_07836_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[16\]
+ net2808 net986 _01309_ VPWR VGND sg13g2_mux2_1
Xhold1767 i_exotiny._0369_\[25\] VPWR VGND net3594 sg13g2_dlygate4sd3_1
X_07767_ net2519 net2780 net990 _01252_ VPWR VGND sg13g2_mux2_1
Xhold1789 i_exotiny.i_wb_spi.dat_rx_r\[27\] VPWR VGND net3616 sg13g2_dlygate4sd3_1
XFILLER_56_267 VPWR VGND sg13g2_fill_2
XFILLER_38_971 VPWR VGND sg13g2_fill_1
X_04979_ VGND VPWR _01424_ _01709_ _01711_ _01388_ sg13g2_a21oi_1
XFILLER_44_407 VPWR VGND sg13g2_fill_2
XFILLER_53_930 VPWR VGND sg13g2_fill_2
X_06718_ net3657 net1102 _02752_ VPWR VGND sg13g2_nor2_1
XFILLER_72_38 VPWR VGND sg13g2_fill_2
XFILLER_24_153 VPWR VGND sg13g2_fill_1
X_07698_ net2172 _03197_ net1000 _01197_ VPWR VGND sg13g2_mux2_1
X_06649_ _01388_ _01467_ _02690_ VPWR VGND sg13g2_nor2_1
XFILLER_24_197 VPWR VGND sg13g2_fill_1
XFILLER_40_668 VPWR VGND sg13g2_fill_2
X_08319_ net359 VGND VPWR net2374 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[21\]
+ clknet_leaf_72_clk_regs sg13g2_dfrbpq_1
X_09299_ net1539 VGND VPWR net2811 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[25\]
+ clknet_leaf_178_clk_regs sg13g2_dfrbpq_1
XFILLER_21_42 VPWR VGND sg13g2_fill_2
XFILLER_106_475 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_102_670 VPWR VGND sg13g2_fill_1
XFILLER_101_191 VPWR VGND sg13g2_decap_8
XFILLER_75_543 VPWR VGND sg13g2_fill_1
XFILLER_75_576 VPWR VGND sg13g2_fill_1
XFILLER_28_481 VPWR VGND sg13g2_fill_2
XFILLER_44_941 VPWR VGND sg13g2_fill_1
XFILLER_71_793 VPWR VGND sg13g2_fill_2
XFILLER_30_134 VPWR VGND sg13g2_fill_2
X_08281__397 VPWR VGND net397 sg13g2_tiehi
XFILLER_8_864 VPWR VGND sg13g2_fill_2
X_08693__1295 VPWR VGND net1715 sg13g2_tiehi
Xhold308 _01297_ VPWR VGND net2135 sg13g2_dlygate4sd3_1
Xhold319 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[4\]
+ VPWR VGND net2146 sg13g2_dlygate4sd3_1
X_08882__1100 VPWR VGND net1520 sg13g2_tiehi
XFILLER_100_629 VPWR VGND sg13g2_fill_1
Xhold1019 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[19\]
+ VPWR VGND net2846 sg13g2_dlygate4sd3_1
X_05951_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[16\]
+ net3283 net970 _00160_ VPWR VGND sg13g2_mux2_1
Xhold1008 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[4\]
+ VPWR VGND net2835 sg13g2_dlygate4sd3_1
X_08670_ net1203 VGND VPWR i_exotiny._2043_\[7\] i_exotiny._2034_\[7\] net1229 sg13g2_dfrbpq_2
X_04902_ net1255 _01613_ _01616_ _01634_ VPWR VGND sg13g2_nor3_2
X_05882_ _02468_ _02431_ _01835_ _01836_ _01496_ VPWR VGND sg13g2_a22oi_1
XFILLER_94_885 VPWR VGND sg13g2_decap_8
X_07621_ _03183_ _03184_ _01133_ VPWR VGND sg13g2_nor2_1
X_04833_ i_exotiny.i_wb_spi.cnt_presc_r\[3\] _01572_ _01573_ VPWR VGND sg13g2_nor2b_1
X_07552_ net3763 _03139_ _03140_ VPWR VGND sg13g2_and2_1
XFILLER_81_535 VPWR VGND sg13g2_fill_1
X_06503_ i_exotiny._0041_\[1\] net883 _02614_ _02617_ VPWR VGND sg13g2_mux2_1
X_04764_ VGND VPWR _01514_ _01515_ net1271 _01369_ sg13g2_a21oi_2
X_08507__173 VPWR VGND net173 sg13g2_tiehi
X_04695_ net1187 _01452_ _01448_ _01453_ VPWR VGND sg13g2_nand3_1
X_07483_ _03108_ VPWR _01071_ VGND _01393_ net903 sg13g2_o21ai_1
X_09222_ net757 VGND VPWR _01277_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[12\]
+ clknet_leaf_136_clk_regs sg13g2_dfrbpq_1
X_06434_ VGND VPWR net1165 _02609_ _02608_ net1138 sg13g2_a21oi_2
X_06365_ net2995 net2493 net1028 _00495_ VPWR VGND sg13g2_mux2_1
X_09153_ net829 VGND VPWR net2546 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[9\]
+ clknet_leaf_172_clk_regs sg13g2_dfrbpq_1
X_08104_ net590 VGND VPWR _00185_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[9\]
+ clknet_leaf_125_clk_regs sg13g2_dfrbpq_1
X_05316_ _01825_ _02039_ _02040_ _02041_ VPWR VGND sg13g2_or3_1
X_06296_ i_exotiny._0016_\[0\] net888 _02552_ _02554_ VPWR VGND sg13g2_mux2_1
X_09084_ net1318 VGND VPWR net2098 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[4\]
+ clknet_leaf_141_clk_regs sg13g2_dfrbpq_1
X_08035_ net659 VGND VPWR _00116_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[4\]
+ clknet_leaf_54_clk_regs sg13g2_dfrbpq_1
Xhold820 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[7\]
+ VPWR VGND net2647 sg13g2_dlygate4sd3_1
X_05247_ net1109 _01969_ _01974_ VPWR VGND sg13g2_and2_1
XFILLER_104_902 VPWR VGND sg13g2_decap_8
Xhold831 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[31\]
+ VPWR VGND net2658 sg13g2_dlygate4sd3_1
Xhold864 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[10\]
+ VPWR VGND net2691 sg13g2_dlygate4sd3_1
Xhold853 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[25\]
+ VPWR VGND net2680 sg13g2_dlygate4sd3_1
X_05178_ _01831_ _01902_ _01903_ _01906_ VPWR VGND sg13g2_nor3_1
Xhold842 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[25\]
+ VPWR VGND net2669 sg13g2_dlygate4sd3_1
XFILLER_103_423 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_93_clk_regs clknet_5_30__leaf_clk_regs clknet_leaf_93_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold886 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[21\]
+ VPWR VGND net2713 sg13g2_dlygate4sd3_1
Xhold897 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[6\]
+ VPWR VGND net2724 sg13g2_dlygate4sd3_1
Xhold875 _00602_ VPWR VGND net2702 sg13g2_dlygate4sd3_1
XFILLER_104_979 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_22_clk_regs clknet_5_12__leaf_clk_regs clknet_leaf_22_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08576__52 VPWR VGND net52 sg13g2_tiehi
X_08514__166 VPWR VGND net166 sg13g2_tiehi
X_08937_ net1465 VGND VPWR net2203 i_exotiny._0042_\[3\] clknet_leaf_52_clk_regs sg13g2_dfrbpq_2
XFILLER_85_830 VPWR VGND sg13g2_fill_1
XFILLER_85_841 VPWR VGND sg13g2_fill_2
X_08868_ net1536 VGND VPWR net3743 i_exotiny.gpo\[1\] clknet_leaf_29_clk_regs sg13g2_dfrbpq_1
Xhold1553 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[16\]
+ VPWR VGND net3380 sg13g2_dlygate4sd3_1
Xhold1531 i_exotiny._0314_\[20\] VPWR VGND net3358 sg13g2_dlygate4sd3_1
Xhold1542 _00828_ VPWR VGND net3369 sg13g2_dlygate4sd3_1
Xhold1520 _00553_ VPWR VGND net3347 sg13g2_dlygate4sd3_1
Xhold1586 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[24\]
+ VPWR VGND net3413 sg13g2_dlygate4sd3_1
Xhold1564 i_exotiny._1465_ VPWR VGND net3391 sg13g2_dlygate4sd3_1
Xhold1575 i_exotiny._0314_\[18\] VPWR VGND net3402 sg13g2_dlygate4sd3_1
X_07819_ net2704 _03220_ net892 _01295_ VPWR VGND sg13g2_mux2_1
Xhold1597 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[21\]
+ VPWR VGND net3424 sg13g2_dlygate4sd3_1
XFILLER_72_524 VPWR VGND sg13g2_fill_2
X_08799_ net1609 VGND VPWR _00857_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[30\]
+ clknet_leaf_163_clk_regs sg13g2_dfrbpq_1
XFILLER_13_657 VPWR VGND sg13g2_fill_2
X_08960__1022 VPWR VGND net1442 sg13g2_tiehi
X_08521__159 VPWR VGND net159 sg13g2_tiehi
XFILLER_5_889 VPWR VGND sg13g2_decap_8
XFILLER_106_272 VPWR VGND sg13g2_decap_8
XFILLER_80_1019 VPWR VGND sg13g2_decap_8
X_08678__1310 VPWR VGND net1730 sg13g2_tiehi
X_08096__598 VPWR VGND net598 sg13g2_tiehi
XFILLER_79_178 VPWR VGND sg13g2_fill_1
XFILLER_29_790 VPWR VGND sg13g2_fill_2
XFILLER_35_248 VPWR VGND sg13g2_fill_1
XFILLER_16_495 VPWR VGND sg13g2_fill_1
X_08780__1208 VPWR VGND net1628 sg13g2_tiehi
X_06150_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[4\] _02476_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[3\]
+ _02533_ VPWR VGND sg13g2_nand3_1
Xhold105 _00061_ VPWR VGND net1932 sg13g2_dlygate4sd3_1
Xhold116 i_exotiny._1924_\[9\] VPWR VGND net1943 sg13g2_dlygate4sd3_1
X_06081_ net2303 net2761 net960 _00257_ VPWR VGND sg13g2_mux2_1
XFILLER_7_193 VPWR VGND sg13g2_fill_1
X_05101_ _01831_ i_exotiny._0550_ _01829_ VPWR VGND sg13g2_nand2_2
Xhold127 _00038_ VPWR VGND net1954 sg13g2_dlygate4sd3_1
Xhold149 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[20\]
+ VPWR VGND net1976 sg13g2_dlygate4sd3_1
Xhold138 i_exotiny._0314_\[26\] VPWR VGND net1965 sg13g2_dlygate4sd3_1
X_05032_ _01764_ i_exotiny._0029_\[3\] _01763_ VPWR VGND sg13g2_nand2_1
XFILLER_99_933 VPWR VGND sg13g2_decap_8
XFILLER_98_432 VPWR VGND sg13g2_decap_8
XFILLER_101_927 VPWR VGND sg13g2_decap_8
X_06983_ net2656 net2742 net1018 _00756_ VPWR VGND sg13g2_mux2_1
XFILLER_100_437 VPWR VGND sg13g2_decap_8
X_05934_ _02486_ net1139 net1167 _02487_ VPWR VGND sg13g2_a21o_1
X_08838__1148 VPWR VGND net1568 sg13g2_tiehi
X_08558__96 VPWR VGND net96 sg13g2_tiehi
X_08722_ net1686 VGND VPWR _00780_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[17\]
+ clknet_leaf_123_clk_regs sg13g2_dfrbpq_1
XFILLER_67_896 VPWR VGND sg13g2_fill_1
XFILLER_96_1026 VPWR VGND sg13g2_fill_2
XFILLER_82_844 VPWR VGND sg13g2_fill_1
XFILLER_82_833 VPWR VGND sg13g2_fill_1
X_08653_ net1744 VGND VPWR _00721_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[22\]
+ clknet_leaf_149_clk_regs sg13g2_dfrbpq_1
X_05865_ _02452_ VPWR _02453_ VGND net3 _01473_ sg13g2_o21ai_1
X_07604_ net1206 net1891 _03173_ _01127_ VPWR VGND sg13g2_nor3_1
X_05796_ _02413_ VPWR _00079_ VGND _00023_ _01551_ sg13g2_o21ai_1
X_04816_ VGND VPWR net1281 i_exotiny._1793_ _01558_ net1265 sg13g2_a21oi_1
X_08584_ net1814 VGND VPWR net2003 i_exotiny._0314_\[29\] clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
XFILLER_82_899 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_140_clk_regs clknet_5_17__leaf_clk_regs clknet_leaf_140_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_22_410 VPWR VGND sg13g2_fill_1
X_04747_ _01471_ _01478_ net1202 _01501_ VPWR VGND _01500_ sg13g2_nand4_1
X_07535_ VGND VPWR _03129_ net3824 net3832 sg13g2_or2_1
X_09286__42 VPWR VGND net42 sg13g2_tiehi
X_07466_ _03099_ _03100_ _03078_ _01062_ VPWR VGND sg13g2_nand3_1
X_09205_ net776 VGND VPWR net2560 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[27\]
+ clknet_leaf_77_clk_regs sg13g2_dfrbpq_1
X_06417_ _02595_ net3551 _02598_ _00515_ VPWR VGND sg13g2_a21o_1
X_04678_ net3523 net3677 net1984 _01439_ VPWR VGND sg13g2_nor3_1
X_08756__1232 VPWR VGND net1652 sg13g2_tiehi
X_07397_ i_exotiny._1160_\[12\] net1216 _03049_ VPWR VGND sg13g2_nor2_1
X_06348_ net3539 i_exotiny._0035_\[3\] net1031 _00478_ VPWR VGND sg13g2_mux2_1
X_09136_ net846 VGND VPWR _01191_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[24\]
+ clknet_leaf_151_clk_regs sg13g2_dfrbpq_1
X_09067_ net1335 VGND VPWR net2030 i_exotiny.i_wdg_top.clk_div_inst.cnt\[7\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_1
X_06279_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[15\]
+ net2385 net942 _00422_ VPWR VGND sg13g2_mux2_1
X_08018_ net676 VGND VPWR net2288 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[19\]
+ clknet_leaf_61_clk_regs sg13g2_dfrbpq_1
Xhold650 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[30\]
+ VPWR VGND net2477 sg13g2_dlygate4sd3_1
Xhold661 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[27\]
+ VPWR VGND net2488 sg13g2_dlygate4sd3_1
Xhold672 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[22\]
+ VPWR VGND net2499 sg13g2_dlygate4sd3_1
XFILLER_103_220 VPWR VGND sg13g2_decap_8
Xhold683 _00142_ VPWR VGND net2510 sg13g2_dlygate4sd3_1
XFILLER_2_859 VPWR VGND sg13g2_decap_8
X_08789__1199 VPWR VGND net1619 sg13g2_tiehi
Xhold694 i_exotiny._0025_\[2\] VPWR VGND net2521 sg13g2_dlygate4sd3_1
XFILLER_104_776 VPWR VGND sg13g2_decap_8
XFILLER_103_297 VPWR VGND sg13g2_decap_8
XFILLER_76_148 VPWR VGND sg13g2_fill_1
X_08978__1004 VPWR VGND net1424 sg13g2_tiehi
XFILLER_92_619 VPWR VGND sg13g2_fill_1
XFILLER_73_800 VPWR VGND sg13g2_fill_2
Xhold1361 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[19\]
+ VPWR VGND net3188 sg13g2_dlygate4sd3_1
XFILLER_57_340 VPWR VGND sg13g2_fill_2
Xhold1350 _01206_ VPWR VGND net3177 sg13g2_dlygate4sd3_1
Xhold1372 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[15\]
+ VPWR VGND net3199 sg13g2_dlygate4sd3_1
Xhold1383 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[6\]
+ VPWR VGND net3210 sg13g2_dlygate4sd3_1
Xhold1394 _01095_ VPWR VGND net3221 sg13g2_dlygate4sd3_1
XFILLER_45_579 VPWR VGND sg13g2_decap_4
XFILLER_72_376 VPWR VGND sg13g2_fill_2
X_08167__511 VPWR VGND net511 sg13g2_tiehi
XFILLER_14_988 VPWR VGND sg13g2_decap_8
X_10675_ i_exotiny.i_wb_spi.sck_r net24 VPWR VGND sg13g2_buf_1
XFILLER_13_487 VPWR VGND sg13g2_fill_2
Xclkbuf_4_6_0_clk_regs clknet_0_clk_regs clknet_4_6_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_96_914 VPWR VGND sg13g2_decap_8
XFILLER_36_502 VPWR VGND sg13g2_fill_1
X_05650_ VGND VPWR net1066 _02307_ _00038_ _02308_ sg13g2_a21oi_1
X_08834__1154 VPWR VGND net1574 sg13g2_tiehi
X_05581_ _01402_ net1204 i_exotiny._2032_ VPWR VGND sg13g2_nor2_1
X_04601_ VPWR _01363_ net3824 VGND sg13g2_inv_1
X_07320_ _02986_ VPWR _01030_ VGND _01382_ net1150 sg13g2_o21ai_1
X_08504__176 VPWR VGND net176 sg13g2_tiehi
X_07251_ net2339 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[14\]
+ net1003 _00974_ VPWR VGND sg13g2_mux2_1
XFILLER_76_0 VPWR VGND sg13g2_fill_2
X_07182_ _02955_ net2106 net1285 VPWR VGND sg13g2_nand2_1
X_06202_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[14\]
+ net2427 net948 _00357_ VPWR VGND sg13g2_mux2_1
XFILLER_9_981 VPWR VGND sg13g2_decap_8
X_06133_ net2709 net3005 net1043 _00302_ VPWR VGND sg13g2_mux2_1
XFILLER_105_529 VPWR VGND sg13g2_decap_8
X_06064_ net2521 net877 _02510_ _02514_ VPWR VGND sg13g2_mux2_1
X_05015_ VGND VPWR _01371_ _01739_ _01747_ _01746_ sg13g2_a21oi_1
XFILLER_101_757 VPWR VGND sg13g2_fill_2
XFILLER_100_234 VPWR VGND sg13g2_decap_8
X_08511__169 VPWR VGND net169 sg13g2_tiehi
X_06966_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[8\]
+ net3099 net1021 _00739_ VPWR VGND sg13g2_mux2_1
XFILLER_104_57 VPWR VGND sg13g2_fill_2
X_05917_ net2123 net2481 net974 _00134_ VPWR VGND sg13g2_mux2_1
X_06897_ _02900_ _02719_ _02462_ net1068 net3817 VPWR VGND sg13g2_a22oi_1
X_08705_ net1703 VGND VPWR net2060 i_exotiny._0032_\[0\] clknet_leaf_120_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_54_354 VPWR VGND sg13g2_fill_1
X_08636_ net1761 VGND VPWR _00704_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[5\]
+ clknet_leaf_147_clk_regs sg13g2_dfrbpq_1
XFILLER_27_557 VPWR VGND sg13g2_fill_2
X_05848_ _02437_ _02433_ _02436_ net1184 _01418_ VPWR VGND sg13g2_a22oi_1
XFILLER_54_365 VPWR VGND sg13g2_decap_4
X_05779_ net3752 VPWR _00072_ VGND net1143 _02402_ sg13g2_o21ai_1
X_08567_ net70 VGND VPWR net3448 i_exotiny._0314_\[12\] clknet_leaf_4_clk_regs sg13g2_dfrbpq_1
X_08498_ net182 VGND VPWR _00572_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[18\]
+ clknet_leaf_93_clk_regs sg13g2_dfrbpq_1
X_07518_ _03114_ VPWR _01098_ VGND _03115_ _03116_ sg13g2_o21ai_1
X_07449_ VGND VPWR net3598 net1083 _03089_ _03077_ sg13g2_a21oi_1
X_09119_ net863 VGND VPWR _01174_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[7\]
+ clknet_leaf_155_clk_regs sg13g2_dfrbpq_1
Xhold480 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[7\]
+ VPWR VGND net2307 sg13g2_dlygate4sd3_1
Xhold491 _00283_ VPWR VGND net2318 sg13g2_dlygate4sd3_1
Xfanout960 _02520_ net960 VPWR VGND sg13g2_buf_8
XFILLER_93_928 VPWR VGND sg13g2_decap_8
Xfanout971 _02487_ net971 VPWR VGND sg13g2_buf_8
XFILLER_77_468 VPWR VGND sg13g2_fill_1
Xfanout982 _03229_ net982 VPWR VGND sg13g2_buf_8
Xfanout993 net994 net993 VPWR VGND sg13g2_buf_8
XFILLER_38_73 VPWR VGND sg13g2_decap_8
Xhold1180 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[28\]
+ VPWR VGND net3007 sg13g2_dlygate4sd3_1
XFILLER_57_192 VPWR VGND sg13g2_fill_1
Xhold1191 _01293_ VPWR VGND net3018 sg13g2_dlygate4sd3_1
XFILLER_73_674 VPWR VGND sg13g2_fill_2
XFILLER_72_162 VPWR VGND sg13g2_fill_1
Xclkload25 clkload25/Y clknet_leaf_45_clk_regs VPWR VGND sg13g2_inv_2
Xclkload14 clkload14/Y clknet_leaf_17_clk_regs VPWR VGND sg13g2_inv_2
XFILLER_10_991 VPWR VGND sg13g2_decap_8
XFILLER_9_299 VPWR VGND sg13g2_fill_2
XFILLER_86_1025 VPWR VGND sg13g2_decap_4
XFILLER_6_962 VPWR VGND sg13g2_decap_8
Xclkload36 VPWR clkload36/Y clknet_leaf_137_clk_regs VGND sg13g2_inv_1
XFILLER_68_424 VPWR VGND sg13g2_fill_2
XFILLER_95_243 VPWR VGND sg13g2_fill_2
X_06820_ VGND VPWR net1097 _02836_ _00679_ _02837_ sg13g2_a21oi_1
X_06751_ net1171 VPWR _02779_ VGND net1933 net1185 sg13g2_o21ai_1
X_05702_ VGND VPWR net1059 _02347_ _00051_ _02345_ sg13g2_a21oi_1
X_06682_ _01506_ _02718_ _02719_ VPWR VGND sg13g2_nor2_2
X_08421_ net264 VGND VPWR _00495_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[20\]
+ clknet_leaf_91_clk_regs sg13g2_dfrbpq_1
X_05633_ VGND VPWR i_exotiny._1615_\[0\] net1125 _02296_ _02295_ sg13g2_a21oi_1
X_08352_ net326 VGND VPWR net3230 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[22\]
+ clknet_leaf_107_clk_regs sg13g2_dfrbpq_1
X_05564_ i_exotiny._0327_\[0\] net1201 _02245_ VPWR VGND sg13g2_nor2_1
X_07303_ net890 i_exotiny._0042_\[0\] _02978_ _02980_ VPWR VGND sg13g2_mux2_1
X_08283_ net395 VGND VPWR _00364_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[17\]
+ clknet_leaf_99_clk_regs sg13g2_dfrbpq_1
X_05495_ _02191_ net3675 net1070 VPWR VGND sg13g2_nand2_1
X_07234_ i_exotiny.i_wb_spi.dat_rx_r\[30\] net3530 net1092 _00959_ VPWR VGND sg13g2_mux2_1
Xclkload8 VPWR clkload8/Y clknet_leaf_180_clk_regs VGND sg13g2_inv_1
X_07165_ net2608 net2052 net1010 _00913_ VPWR VGND sg13g2_mux2_1
XFILLER_105_326 VPWR VGND sg13g2_decap_8
X_06116_ net2115 i_exotiny._0037_\[3\] net1046 _00285_ VPWR VGND sg13g2_mux2_1
X_07096_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[24\]
+ net2694 net914 _00851_ VPWR VGND sg13g2_mux2_1
X_08157__521 VPWR VGND net521 sg13g2_tiehi
X_06047_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[19\]
+ net3060 net963 _00232_ VPWR VGND sg13g2_mux2_1
XFILLER_8_1014 VPWR VGND sg13g2_decap_8
X_07998_ i_exotiny._2032_ VGND VPWR i_exotiny._2044_\[1\] i_exotiny.i_wdg_top.cntr_inst.rst_n_sync
+ net1228 sg13g2_dfrbpq_2
X_06949_ net2734 _02918_ net926 _00727_ VPWR VGND sg13g2_mux2_1
X_08619_ net1777 VGND VPWR net3748 i_exotiny._1619_\[3\] clknet_leaf_21_clk_regs sg13g2_dfrbpq_2
XFILLER_30_519 VPWR VGND sg13g2_decap_4
X_08164__514 VPWR VGND net514 sg13g2_tiehi
XFILLER_23_582 VPWR VGND sg13g2_fill_1
XFILLER_10_243 VPWR VGND sg13g2_fill_1
XFILLER_10_254 VPWR VGND sg13g2_fill_2
XFILLER_40_30 VPWR VGND sg13g2_fill_2
XFILLER_40_41 VPWR VGND sg13g2_fill_2
XFILLER_3_921 VPWR VGND sg13g2_decap_8
X_09270__81 VPWR VGND net81 sg13g2_tiehi
XFILLER_105_860 VPWR VGND sg13g2_decap_8
XFILLER_3_998 VPWR VGND sg13g2_decap_8
XFILLER_78_755 VPWR VGND sg13g2_fill_1
XFILLER_93_703 VPWR VGND sg13g2_fill_1
XFILLER_77_298 VPWR VGND sg13g2_fill_2
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_53_1002 VPWR VGND sg13g2_fill_2
X_08540__140 VPWR VGND net140 sg13g2_tiehi
XFILLER_14_1019 VPWR VGND sg13g2_decap_8
X_08501__179 VPWR VGND net179 sg13g2_tiehi
X_05280_ _02006_ _01784_ i_exotiny._0042_\[0\] _01771_ i_exotiny._0016_\[0\] VPWR
+ VGND sg13g2_a22oi_1
Xclkbuf_5_2__f_clk_regs clknet_4_1_0_clk_regs clknet_5_2__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08970_ net1432 VGND VPWR net3685 i_exotiny._0590_ clknet_leaf_12_clk_regs sg13g2_dfrbpq_2
XFILLER_102_329 VPWR VGND sg13g2_decap_8
X_07921_ net727 VGND VPWR net1940 i_exotiny._1924_\[14\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
XFILLER_96_563 VPWR VGND sg13g2_fill_2
Xhold1905 i_exotiny._1652_\[0\] VPWR VGND net3732 sg13g2_dlygate4sd3_1
Xhold1916 _00926_ VPWR VGND net3743 sg13g2_dlygate4sd3_1
XFILLER_29_608 VPWR VGND sg13g2_fill_1
X_07852_ i_exotiny._0022_\[0\] net889 _03222_ _03224_ VPWR VGND sg13g2_mux2_1
Xhold1927 i_exotiny._1309_ VPWR VGND net3754 sg13g2_dlygate4sd3_1
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_1
X_06803_ VGND VPWR _01417_ net1191 _02823_ _01517_ sg13g2_a21oi_1
XFILLER_56_427 VPWR VGND sg13g2_decap_4
Xhold1938 _00509_ VPWR VGND net3765 sg13g2_dlygate4sd3_1
Xhold1949 _02605_ VPWR VGND net3776 sg13g2_dlygate4sd3_1
X_07783_ _03215_ net2853 net988 _01264_ VPWR VGND sg13g2_mux2_1
XFILLER_37_641 VPWR VGND sg13g2_decap_4
X_04995_ _01725_ _01726_ _01711_ _01727_ VPWR VGND sg13g2_nand3_1
XFILLER_65_983 VPWR VGND sg13g2_fill_1
X_06734_ VGND VPWR net1980 net1137 _02765_ _02764_ sg13g2_a21oi_1
XFILLER_80_931 VPWR VGND sg13g2_fill_1
X_06665_ _02691_ VPWR _02704_ VGND _02688_ _02702_ sg13g2_o21ai_1
XFILLER_36_184 VPWR VGND sg13g2_fill_1
X_08404_ net281 VGND VPWR net3540 i_exotiny._0035_\[3\] clknet_leaf_96_clk_regs sg13g2_dfrbpq_2
X_05616_ net1120 net1907 _02283_ VPWR VGND sg13g2_nor2b_1
XFILLER_52_688 VPWR VGND sg13g2_fill_2
XFILLER_12_508 VPWR VGND sg13g2_fill_2
X_08335_ net343 VGND VPWR _00416_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[5\]
+ clknet_leaf_108_clk_regs sg13g2_dfrbpq_1
X_06596_ net3498 net1155 _02654_ VPWR VGND sg13g2_nor2_1
X_05547_ _02231_ VPWR _02232_ VGND net1275 i_exotiny._0315_\[19\] sg13g2_o21ai_1
X_08266_ net412 VGND VPWR net2147 i_exotiny._0033_\[0\] clknet_leaf_101_clk_regs sg13g2_dfrbpq_2
X_05478_ net3707 _02177_ _02179_ VPWR VGND sg13g2_nor2_1
X_07217_ VGND VPWR _01416_ net1090 _00944_ _02969_ sg13g2_a21oi_1
X_08197_ net480 VGND VPWR _00278_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[28\]
+ clknet_leaf_110_clk_regs sg13g2_dfrbpq_1
X_07148_ net2828 net2204 net1012 _00896_ VPWR VGND sg13g2_mux2_1
XFILLER_106_657 VPWR VGND sg13g2_decap_8
XFILLER_105_123 VPWR VGND sg13g2_decap_8
XFILLER_10_44 VPWR VGND sg13g2_fill_1
X_07079_ net2359 net2644 net915 _00834_ VPWR VGND sg13g2_mux2_1
Xfanout1029 net1032 net1029 VPWR VGND sg13g2_buf_8
Xfanout1007 _02973_ net1007 VPWR VGND sg13g2_buf_8
Xfanout1018 net1019 net1018 VPWR VGND sg13g2_buf_8
XFILLER_0_924 VPWR VGND sg13g2_decap_8
XFILLER_102_874 VPWR VGND sg13g2_decap_8
XFILLER_87_541 VPWR VGND sg13g2_decap_4
XFILLER_101_373 VPWR VGND sg13g2_decap_8
XFILLER_87_596 VPWR VGND sg13g2_fill_1
XFILLER_59_298 VPWR VGND sg13g2_fill_2
X_09200__781 VPWR VGND net781 sg13g2_tiehi
XFILLER_43_611 VPWR VGND sg13g2_fill_2
XFILLER_15_324 VPWR VGND sg13g2_fill_1
XFILLER_15_357 VPWR VGND sg13g2_fill_1
XFILLER_43_655 VPWR VGND sg13g2_fill_1
XFILLER_43_699 VPWR VGND sg13g2_decap_8
XFILLER_100_1022 VPWR VGND sg13g2_decap_8
XFILLER_98_839 VPWR VGND sg13g2_decap_8
XFILLER_83_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_250 VPWR VGND sg13g2_fill_2
XFILLER_97_338 VPWR VGND sg13g2_decap_8
XFILLER_3_795 VPWR VGND sg13g2_decap_8
XFILLER_2_283 VPWR VGND sg13g2_fill_1
X_07993__134 VPWR VGND net134 sg13g2_tiehi
XFILLER_19_641 VPWR VGND sg13g2_fill_1
X_04780_ VGND VPWR net1246 _01387_ _01530_ net1273 sg13g2_a21oi_1
XFILLER_61_463 VPWR VGND sg13g2_fill_2
X_06450_ net2679 net2206 net935 _00537_ VPWR VGND sg13g2_mux2_1
X_05401_ i_exotiny._2034_\[4\] _02113_ _02116_ VPWR VGND sg13g2_nor2_1
XFILLER_21_316 VPWR VGND sg13g2_fill_2
XFILLER_22_828 VPWR VGND sg13g2_fill_1
X_08147__531 VPWR VGND net531 sg13g2_tiehi
XFILLER_34_699 VPWR VGND sg13g2_fill_1
X_06381_ _01513_ VPWR _02571_ VGND _01489_ _01521_ sg13g2_o21ai_1
X_05332_ _01388_ VPWR _02056_ VGND i_exotiny._0352_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r
+ sg13g2_o21ai_1
X_08120_ net574 VGND VPWR _00201_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[25\]
+ clknet_leaf_124_clk_regs sg13g2_dfrbpq_1
X_08051_ net643 VGND VPWR _00132_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[20\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
X_05263_ _01989_ i_exotiny._0015_\[0\] _01761_ VPWR VGND sg13g2_nand2_1
X_07002_ net2627 net3178 net919 _00769_ VPWR VGND sg13g2_mux2_1
XFILLER_89_806 VPWR VGND sg13g2_fill_2
X_08914__1068 VPWR VGND net1488 sg13g2_tiehi
Xclkbuf_leaf_165_clk_regs clknet_5_6__leaf_clk_regs clknet_leaf_165_clk_regs VPWR
+ VGND sg13g2_buf_8
X_05194_ _01922_ _01777_ i_exotiny._0013_\[1\] _01770_ i_exotiny._0025_\[1\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_103_649 VPWR VGND sg13g2_decap_4
XFILLER_103_638 VPWR VGND sg13g2_fill_2
X_08953_ net1449 VGND VPWR net2847 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[19\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
XFILLER_102_159 VPWR VGND sg13g2_fill_1
Xhold1702 _00069_ VPWR VGND net3529 sg13g2_dlygate4sd3_1
X_08154__524 VPWR VGND net524 sg13g2_tiehi
X_07904_ net43 VGND VPWR net3696 i_exotiny._1311_ clknet_leaf_6_clk_regs sg13g2_dfrbpq_2
XFILLER_99_1024 VPWR VGND sg13g2_decap_4
XFILLER_96_371 VPWR VGND sg13g2_decap_8
Xhold1713 _00478_ VPWR VGND net3540 sg13g2_dlygate4sd3_1
X_08884_ net1518 VGND VPWR net1946 i_exotiny.i_wb_spi.dat_rx_r\[14\] clknet_leaf_59_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_69_574 VPWR VGND sg13g2_fill_1
Xhold1735 i_exotiny._1902_\[5\] VPWR VGND net3562 sg13g2_dlygate4sd3_1
Xhold1724 i_exotiny._2025_\[3\] VPWR VGND net3551 sg13g2_dlygate4sd3_1
Xhold1746 _00685_ VPWR VGND net3573 sg13g2_dlygate4sd3_1
Xhold1768 i_exotiny._1611_\[5\] VPWR VGND net3595 sg13g2_dlygate4sd3_1
Xhold1757 i_exotiny._0369_\[27\] VPWR VGND net3584 sg13g2_dlygate4sd3_1
X_07835_ net3222 net3137 net983 _01308_ VPWR VGND sg13g2_mux2_1
X_07945__89 VPWR VGND net89 sg13g2_tiehi
X_07766_ net3317 net2581 net989 _01251_ VPWR VGND sg13g2_mux2_1
Xhold1779 i_exotiny._1956_ VPWR VGND net3606 sg13g2_dlygate4sd3_1
X_04978_ VGND VPWR _01710_ _01708_ net1180 sg13g2_or2_1
X_06717_ VGND VPWR net3611 net1137 _02751_ _02750_ sg13g2_a21oi_1
X_07697_ net2511 net877 _03193_ _03197_ VPWR VGND sg13g2_mux2_1
X_06648_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r[0] i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[0\].i_hadd.a_i
+ _02689_ VPWR VGND sg13g2_xor2_1
X_06579_ net1199 _02641_ _02642_ _00633_ VPWR VGND sg13g2_nor3_1
X_08318_ net360 VGND VPWR net2201 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[20\]
+ clknet_leaf_82_clk_regs sg13g2_dfrbpq_1
X_09298_ net1767 VGND VPWR net2254 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[24\]
+ clknet_leaf_178_clk_regs sg13g2_dfrbpq_1
X_08161__517 VPWR VGND net517 sg13g2_tiehi
X_08249_ net428 VGND VPWR net2110 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[16\]
+ clknet_leaf_56_clk_regs sg13g2_dfrbpq_1
XFILLER_20_382 VPWR VGND sg13g2_fill_2
XFILLER_106_454 VPWR VGND sg13g2_decap_8
X_07977__118 VPWR VGND net118 sg13g2_tiehi
XFILLER_0_721 VPWR VGND sg13g2_decap_8
XFILLER_43_1001 VPWR VGND sg13g2_fill_1
XFILLER_102_660 VPWR VGND sg13g2_fill_1
XFILLER_94_319 VPWR VGND sg13g2_decap_8
X_08530__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_35_408 VPWR VGND sg13g2_fill_1
XFILLER_16_677 VPWR VGND sg13g2_fill_1
XFILLER_30_124 VPWR VGND sg13g2_fill_2
Xhold309 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[7\]
+ VPWR VGND net2136 sg13g2_dlygate4sd3_1
XFILLER_3_570 VPWR VGND sg13g2_fill_2
X_05950_ net2822 net2892 net969 _00159_ VPWR VGND sg13g2_mux2_1
Xhold1009 _00590_ VPWR VGND net2836 sg13g2_dlygate4sd3_1
X_05881_ VGND VPWR _01836_ _02269_ _02467_ _02428_ sg13g2_a21oi_1
X_04901_ _01633_ _01632_ i_exotiny._0022_\[3\] _01631_ i_exotiny._0027_\[3\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_93_341 VPWR VGND sg13g2_fill_1
X_07620_ i_exotiny._0000_ VPWR _03184_ VGND net3569 _03182_ sg13g2_o21ai_1
X_04832_ net1840 net3728 net3814 _01572_ VPWR VGND sg13g2_nor3_1
XFILLER_53_205 VPWR VGND sg13g2_fill_2
X_07551_ _03133_ _03138_ _03139_ _01108_ VPWR VGND sg13g2_nor3_1
XFILLER_19_482 VPWR VGND sg13g2_fill_2
X_06502_ _02616_ net2561 net1024 _00582_ VPWR VGND sg13g2_mux2_1
X_04763_ net1272 i_exotiny._0315_\[31\] _01514_ VPWR VGND sg13g2_nor2_1
X_04694_ net3705 net3841 _01452_ VPWR VGND sg13g2_nor2_1
X_07482_ _03108_ net1234 net903 VPWR VGND sg13g2_nand2_1
X_06433_ _02509_ _02518_ _02608_ VPWR VGND sg13g2_nor2_2
X_09221_ net758 VGND VPWR net2252 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[11\]
+ clknet_leaf_137_clk_regs sg13g2_dfrbpq_1
X_06364_ net2515 net2942 net1030 _00494_ VPWR VGND sg13g2_mux2_1
X_09152_ net830 VGND VPWR net2336 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[8\]
+ clknet_leaf_175_clk_regs sg13g2_dfrbpq_1
X_08103_ net591 VGND VPWR net2155 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[8\]
+ clknet_leaf_125_clk_regs sg13g2_dfrbpq_1
X_05315_ _02039_ _02040_ net34 VPWR VGND sg13g2_nor2_2
X_06295_ net2673 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[27\]
+ net942 _00438_ VPWR VGND sg13g2_mux2_1
X_09083_ net1319 VGND VPWR net2918 i_exotiny._0024_\[3\] clknet_leaf_144_clk_regs
+ sg13g2_dfrbpq_2
X_08034_ net660 VGND VPWR net2896 i_exotiny._0019_\[3\] clknet_leaf_54_clk_regs sg13g2_dfrbpq_2
Xhold821 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[18\]
+ VPWR VGND net2648 sg13g2_dlygate4sd3_1
Xhold810 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[4\]
+ VPWR VGND net2637 sg13g2_dlygate4sd3_1
X_05246_ _01973_ net35 _01825_ VPWR VGND sg13g2_nand2b_1
Xhold832 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[26\]
+ VPWR VGND net2659 sg13g2_dlygate4sd3_1
Xhold854 _01290_ VPWR VGND net2681 sg13g2_dlygate4sd3_1
X_05177_ _01831_ VPWR _01905_ VGND _01902_ _01903_ sg13g2_o21ai_1
Xhold843 _00197_ VPWR VGND net2670 sg13g2_dlygate4sd3_1
XFILLER_104_958 VPWR VGND sg13g2_decap_8
XFILLER_103_402 VPWR VGND sg13g2_decap_8
Xhold876 i_exotiny._0041_\[0\] VPWR VGND net2703 sg13g2_dlygate4sd3_1
Xhold887 _00981_ VPWR VGND net2714 sg13g2_dlygate4sd3_1
Xhold898 _01205_ VPWR VGND net2725 sg13g2_dlygate4sd3_1
Xhold865 _00292_ VPWR VGND net2692 sg13g2_dlygate4sd3_1
X_07956__703 VPWR VGND net703 sg13g2_tiehi
XFILLER_103_479 VPWR VGND sg13g2_decap_8
X_08936_ net1466 VGND VPWR _00994_ i_exotiny._0042_\[2\] clknet_leaf_74_clk_regs sg13g2_dfrbpq_2
Xhold1510 i_exotiny._0033_\[2\] VPWR VGND net3337 sg13g2_dlygate4sd3_1
Xhold1543 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[29\]
+ VPWR VGND net3370 sg13g2_dlygate4sd3_1
Xhold1521 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[10\]
+ VPWR VGND net3348 sg13g2_dlygate4sd3_1
X_08867_ net1538 VGND VPWR net3774 i_exotiny.gpo\[0\] clknet_leaf_29_clk_regs sg13g2_dfrbpq_1
Xhold1532 _00644_ VPWR VGND net3359 sg13g2_dlygate4sd3_1
Xhold1565 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[16\]
+ VPWR VGND net3392 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_62_clk_regs clknet_5_13__leaf_clk_regs clknet_leaf_62_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold1554 _00711_ VPWR VGND net3381 sg13g2_dlygate4sd3_1
Xhold1576 _00642_ VPWR VGND net3403 sg13g2_dlygate4sd3_1
X_07818_ i_exotiny._0023_\[2\] net879 _03216_ _03220_ VPWR VGND sg13g2_mux2_1
Xhold1598 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[23\]
+ VPWR VGND net3425 sg13g2_dlygate4sd3_1
Xhold1587 _00847_ VPWR VGND net3414 sg13g2_dlygate4sd3_1
X_08798_ net1610 VGND VPWR net2937 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[29\]
+ clknet_leaf_169_clk_regs sg13g2_dfrbpq_1
X_07749_ net2600 i_exotiny._0026_\[1\] net989 _01234_ VPWR VGND sg13g2_mux2_1
XFILLER_25_485 VPWR VGND sg13g2_fill_2
XFILLER_106_251 VPWR VGND sg13g2_decap_8
XFILLER_106_0 VPWR VGND sg13g2_fill_2
XFILLER_5_868 VPWR VGND sg13g2_decap_8
XFILLER_102_490 VPWR VGND sg13g2_decap_8
XFILLER_29_780 VPWR VGND sg13g2_fill_1
XFILLER_35_216 VPWR VGND sg13g2_fill_2
XFILLER_35_227 VPWR VGND sg13g2_fill_2
XFILLER_48_599 VPWR VGND sg13g2_decap_4
XFILLER_32_967 VPWR VGND sg13g2_fill_2
XFILLER_85_5 VPWR VGND sg13g2_fill_2
XFILLER_89_1023 VPWR VGND sg13g2_decap_4
Xhold117 _00034_ VPWR VGND net1944 sg13g2_dlygate4sd3_1
X_06080_ net2255 net2843 net958 _00256_ VPWR VGND sg13g2_mux2_1
Xhold106 i_exotiny.i_wb_spi.dat_rx_r\[9\] VPWR VGND net1933 sg13g2_dlygate4sd3_1
X_05100_ i_exotiny._0550_ _01829_ _01830_ VPWR VGND sg13g2_and2_1
XFILLER_99_912 VPWR VGND sg13g2_decap_8
Xhold139 _00650_ VPWR VGND net1966 sg13g2_dlygate4sd3_1
X_05031_ net1220 _01759_ _01762_ _01763_ VPWR VGND sg13g2_nor3_2
Xhold128 i_exotiny._1160_\[7\] VPWR VGND net1955 sg13g2_dlygate4sd3_1
XFILLER_98_411 VPWR VGND sg13g2_decap_8
XFILLER_101_906 VPWR VGND sg13g2_decap_8
XFILLER_99_989 VPWR VGND sg13g2_decap_8
XFILLER_4_890 VPWR VGND sg13g2_decap_8
XFILLER_100_416 VPWR VGND sg13g2_decap_8
XFILLER_98_488 VPWR VGND sg13g2_decap_8
X_06982_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[24\]
+ net2355 net1021 _00755_ VPWR VGND sg13g2_mux2_1
XFILLER_66_330 VPWR VGND sg13g2_fill_2
X_05933_ _02477_ _02485_ _02486_ VPWR VGND sg13g2_nor2_2
X_08846__1140 VPWR VGND net1560 sg13g2_tiehi
X_09294__1391 VPWR VGND net1811 sg13g2_tiehi
X_08151__527 VPWR VGND net527 sg13g2_tiehi
X_08721_ net1687 VGND VPWR net2646 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[16\]
+ clknet_leaf_119_clk_regs sg13g2_dfrbpq_1
XFILLER_96_1005 VPWR VGND sg13g2_decap_8
Xfanout1190 net1191 net1190 VPWR VGND sg13g2_buf_8
X_08652_ net1745 VGND VPWR _00720_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[21\]
+ clknet_leaf_148_clk_regs sg13g2_dfrbpq_1
X_07603_ _03173_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[11\] net1890 _03170_ VPWR VGND
+ sg13g2_and3_1
XFILLER_54_536 VPWR VGND sg13g2_fill_1
X_05864_ net1184 _02447_ _02451_ _02452_ VPWR VGND sg13g2_or3_1
X_05795_ _02413_ net1873 net1145 VPWR VGND sg13g2_nand2_1
X_04815_ i_exotiny._1725_ net1264 _01557_ VPWR VGND sg13g2_nor2_1
X_08583_ net1816 VGND VPWR net2447 i_exotiny._0314_\[28\] clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
XFILLER_81_377 VPWR VGND sg13g2_fill_2
XFILLER_22_400 VPWR VGND sg13g2_fill_1
X_04746_ net1224 _01497_ _01500_ VPWR VGND net1254 sg13g2_nand3b_1
X_07534_ VGND VPWR _03127_ _03128_ _01102_ net1196 sg13g2_a21oi_1
X_07465_ _03100_ net1148 _03037_ VPWR VGND sg13g2_nand2_1
X_09204_ net777 VGND VPWR _01259_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[26\]
+ clknet_leaf_76_clk_regs sg13g2_dfrbpq_1
X_06416_ net1282 VPWR _02598_ VGND _01361_ _02595_ sg13g2_o21ai_1
X_04677_ _01438_ _01435_ net3790 _01426_ _01424_ VPWR VGND sg13g2_a22oi_1
X_08520__160 VPWR VGND net160 sg13g2_tiehi
Xclkbuf_leaf_180_clk_regs clknet_5_1__leaf_clk_regs clknet_leaf_180_clk_regs VPWR
+ VGND sg13g2_buf_8
X_07396_ VGND VPWR net1077 _03048_ _01044_ _03043_ sg13g2_a21oi_1
X_06347_ net3373 net3343 net1030 _00477_ VPWR VGND sg13g2_mux2_1
X_09135_ net847 VGND VPWR _01190_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[23\]
+ clknet_leaf_156_clk_regs sg13g2_dfrbpq_1
X_09066_ net1336 VGND VPWR net1915 i_exotiny.i_wdg_top.clk_div_inst.cnt\[6\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_1
X_06278_ net2775 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[10\]
+ net941 _00421_ VPWR VGND sg13g2_mux2_1
X_08017_ net677 VGND VPWR _00098_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[18\]
+ clknet_leaf_61_clk_regs sg13g2_dfrbpq_1
X_05229_ _01957_ _01956_ _01643_ _01650_ i_exotiny._0016_\[1\] VPWR VGND sg13g2_a22oi_1
Xhold651 _00174_ VPWR VGND net2478 sg13g2_dlygate4sd3_1
Xhold662 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[21\]
+ VPWR VGND net2489 sg13g2_dlygate4sd3_1
Xhold640 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[7\]
+ VPWR VGND net2467 sg13g2_dlygate4sd3_1
XFILLER_2_838 VPWR VGND sg13g2_decap_8
XFILLER_104_755 VPWR VGND sg13g2_decap_8
Xhold695 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[31\]
+ VPWR VGND net2522 sg13g2_dlygate4sd3_1
X_08651__1326 VPWR VGND net1746 sg13g2_tiehi
X_08797__1191 VPWR VGND net1611 sg13g2_tiehi
Xhold673 _01189_ VPWR VGND net2500 sg13g2_dlygate4sd3_1
Xhold684 i_exotiny._0030_\[2\] VPWR VGND net2511 sg13g2_dlygate4sd3_1
XFILLER_103_276 VPWR VGND sg13g2_decap_8
XFILLER_89_499 VPWR VGND sg13g2_fill_2
XFILLER_58_853 VPWR VGND sg13g2_fill_1
X_08919_ net1483 VGND VPWR _00977_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[17\]
+ clknet_leaf_113_clk_regs sg13g2_dfrbpq_1
XFILLER_58_864 VPWR VGND sg13g2_fill_1
Xhold1340 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[20\]
+ VPWR VGND net3167 sg13g2_dlygate4sd3_1
XFILLER_40_1026 VPWR VGND sg13g2_fill_2
Xhold1351 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[10\]
+ VPWR VGND net3178 sg13g2_dlygate4sd3_1
XFILLER_100_994 VPWR VGND sg13g2_decap_8
Xhold1373 _00810_ VPWR VGND net3200 sg13g2_dlygate4sd3_1
Xhold1384 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[13\]
+ VPWR VGND net3211 sg13g2_dlygate4sd3_1
XFILLER_73_845 VPWR VGND sg13g2_fill_2
Xhold1362 _00362_ VPWR VGND net3189 sg13g2_dlygate4sd3_1
Xhold1395 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[15\]
+ VPWR VGND net3222 sg13g2_dlygate4sd3_1
X_08873__1109 VPWR VGND net1529 sg13g2_tiehi
XFILLER_14_967 VPWR VGND sg13g2_decap_8
XFILLER_25_293 VPWR VGND sg13g2_fill_1
XFILLER_41_742 VPWR VGND sg13g2_fill_2
X_10674_ ccx_req net23 VPWR VGND sg13g2_buf_1
XFILLER_95_414 VPWR VGND sg13g2_fill_2
XFILLER_49_886 VPWR VGND sg13g2_fill_1
XFILLER_76_694 VPWR VGND sg13g2_fill_2
XFILLER_36_536 VPWR VGND sg13g2_fill_2
XFILLER_1_1020 VPWR VGND sg13g2_decap_8
XFILLER_63_377 VPWR VGND sg13g2_fill_2
X_04600_ _01362_ net3834 VPWR VGND sg13g2_inv_2
X_05580_ i_exotiny._1793_ net1218 _01555_ _10677_/A VPWR VGND sg13g2_or3_1
XFILLER_17_1017 VPWR VGND sg13g2_fill_2
X_07250_ net2924 net3089 net1005 _00973_ VPWR VGND sg13g2_mux2_1
XFILLER_20_948 VPWR VGND sg13g2_fill_1
X_06201_ net3186 net2947 net946 _00356_ VPWR VGND sg13g2_mux2_1
X_07181_ net3622 net3656 _02954_ _00923_ VPWR VGND sg13g2_mux2_1
XFILLER_9_960 VPWR VGND sg13g2_decap_8
XFILLER_69_0 VPWR VGND sg13g2_fill_2
X_06132_ net3503 net3454 net1044 _00301_ VPWR VGND sg13g2_mux2_1
XFILLER_105_508 VPWR VGND sg13g2_decap_8
X_06063_ _02513_ net2795 net962 _00246_ VPWR VGND sg13g2_mux2_1
X_05014_ _01746_ _01425_ _01710_ VPWR VGND sg13g2_nand2_1
XFILLER_63_1026 VPWR VGND sg13g2_fill_2
XFILLER_98_285 VPWR VGND sg13g2_decap_8
X_06965_ net3247 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[11\]
+ net1019 _00738_ VPWR VGND sg13g2_mux2_1
X_08704_ net1704 VGND VPWR _00762_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[31\]
+ clknet_leaf_105_clk_regs sg13g2_dfrbpq_1
XFILLER_104_69 VPWR VGND sg13g2_fill_2
X_05916_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[21\]
+ net2164 net972 _00133_ VPWR VGND sg13g2_mux2_1
X_06896_ _02899_ VPWR _00693_ VGND _02453_ _02720_ sg13g2_o21ai_1
XFILLER_27_536 VPWR VGND sg13g2_fill_2
XFILLER_39_363 VPWR VGND sg13g2_fill_1
X_08635_ net1762 VGND VPWR _00703_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[4\]
+ clknet_leaf_143_clk_regs sg13g2_dfrbpq_1
X_05847_ VGND VPWR _02434_ _02435_ _02436_ net1184 sg13g2_a21oi_1
X_08566_ net72 VGND VPWR net3499 i_exotiny._0314_\[11\] clknet_leaf_179_clk_regs sg13g2_dfrbpq_2
X_05778_ _02403_ net1126 _01375_ net1145 net3751 VPWR VGND sg13g2_a22oi_1
X_07517_ _03106_ VPWR _03116_ VGND _01500_ _02014_ sg13g2_o21ai_1
X_08497_ net183 VGND VPWR _00571_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[17\]
+ clknet_leaf_71_clk_regs sg13g2_dfrbpq_1
X_04729_ _01485_ net3754 _01464_ VPWR VGND sg13g2_nand2_2
XFILLER_50_594 VPWR VGND sg13g2_fill_1
XFILLER_50_572 VPWR VGND sg13g2_fill_1
X_07448_ _03088_ net1149 _03021_ net1209 net3384 VPWR VGND sg13g2_a22oi_1
XFILLER_10_436 VPWR VGND sg13g2_fill_2
XFILLER_7_919 VPWR VGND sg13g2_decap_8
X_08705__1283 VPWR VGND net1703 sg13g2_tiehi
X_07379_ i_exotiny._0369_\[28\] net1213 _03035_ VPWR VGND sg13g2_and2_1
X_09118_ net864 VGND VPWR _01173_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[6\]
+ clknet_leaf_156_clk_regs sg13g2_dfrbpq_1
X_09049_ net1354 VGND VPWR i_exotiny._1266_ i_exotiny._0352_ clknet_leaf_4_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_104_530 VPWR VGND sg13g2_decap_8
X_08600__1376 VPWR VGND net1796 sg13g2_tiehi
Xhold470 _01165_ VPWR VGND net2297 sg13g2_dlygate4sd3_1
Xhold481 _01300_ VPWR VGND net2308 sg13g2_dlygate4sd3_1
XFILLER_104_563 VPWR VGND sg13g2_decap_8
Xhold492 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[8\]
+ VPWR VGND net2319 sg13g2_dlygate4sd3_1
Xfanout950 net951 net950 VPWR VGND sg13g2_buf_8
Xfanout961 net965 net961 VPWR VGND sg13g2_buf_8
Xfanout972 net977 net972 VPWR VGND sg13g2_buf_8
X_08927__1055 VPWR VGND net1475 sg13g2_tiehi
Xfanout994 net997 net994 VPWR VGND sg13g2_buf_8
Xfanout983 net985 net983 VPWR VGND sg13g2_buf_8
Xhold1170 i_exotiny._0369_\[9\] VPWR VGND net2997 sg13g2_dlygate4sd3_1
XFILLER_38_96 VPWR VGND sg13g2_fill_1
Xhold1181 _01261_ VPWR VGND net3008 sg13g2_dlygate4sd3_1
Xhold1192 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[9\]
+ VPWR VGND net3019 sg13g2_dlygate4sd3_1
XFILLER_57_182 VPWR VGND sg13g2_decap_4
XFILLER_46_856 VPWR VGND sg13g2_fill_1
XFILLER_60_336 VPWR VGND sg13g2_fill_1
X_08386__292 VPWR VGND net292 sg13g2_tiehi
XFILLER_70_50 VPWR VGND sg13g2_fill_2
XFILLER_70_72 VPWR VGND sg13g2_fill_2
Xclkload26 clkload26/Y clknet_leaf_21_clk_regs VPWR VGND sg13g2_inv_2
XFILLER_10_970 VPWR VGND sg13g2_decap_8
Xclkload15 clkload15/Y clknet_leaf_162_clk_regs VPWR VGND sg13g2_inv_2
XFILLER_86_1004 VPWR VGND sg13g2_decap_8
Xclkload37 VPWR clkload37/Y clknet_leaf_104_clk_regs VGND sg13g2_inv_1
XFILLER_6_941 VPWR VGND sg13g2_decap_8
Xclkbuf_5_1__f_clk_regs clknet_4_0_0_clk_regs clknet_5_1__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_5_495 VPWR VGND sg13g2_fill_1
XFILLER_95_233 VPWR VGND sg13g2_fill_1
X_08510__170 VPWR VGND net170 sg13g2_tiehi
X_06750_ VGND VPWR net1100 _02777_ _00668_ _02778_ sg13g2_a21oi_1
XFILLER_55_119 VPWR VGND sg13g2_fill_1
XFILLER_55_108 VPWR VGND sg13g2_fill_2
XFILLER_49_672 VPWR VGND sg13g2_decap_4
XFILLER_36_300 VPWR VGND sg13g2_fill_1
X_05701_ VGND VPWR i_exotiny._1619_\[1\] net1117 _02347_ _02346_ sg13g2_a21oi_1
Xclkbuf_leaf_119_clk_regs clknet_5_20__leaf_clk_regs clknet_leaf_119_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_37_867 VPWR VGND sg13g2_fill_1
X_06681_ _02718_ net1102 VPWR VGND sg13g2_inv_2
XFILLER_93_1019 VPWR VGND sg13g2_decap_8
XFILLER_92_984 VPWR VGND sg13g2_decap_8
X_05632_ net1124 net1941 _02295_ VPWR VGND sg13g2_nor2b_1
X_08420_ net265 VGND VPWR _00494_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[19\]
+ clknet_leaf_97_clk_regs sg13g2_dfrbpq_1
X_08351_ net327 VGND VPWR net2368 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[21\]
+ clknet_leaf_94_clk_regs sg13g2_dfrbpq_1
X_05563_ _02244_ i_exotiny._0315_\[7\] _01690_ VPWR VGND sg13g2_xnor2_1
X_07302_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[27\]
+ net2495 net911 _01019_ VPWR VGND sg13g2_mux2_1
X_08282_ net396 VGND VPWR _00363_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[16\]
+ clknet_leaf_100_clk_regs sg13g2_dfrbpq_1
XFILLER_20_712 VPWR VGND sg13g2_fill_2
X_05494_ _02188_ VPWR i_exotiny._1611_\[11\] VGND net1075 _02190_ sg13g2_o21ai_1
X_07233_ i_exotiny.i_wb_spi.dat_rx_r\[29\] net3582 net1092 _00958_ VPWR VGND sg13g2_mux2_1
Xclkload9 clkload9/Y clknet_leaf_4_clk_regs VPWR VGND sg13g2_inv_2
X_07164_ net3160 net2213 net1008 _00912_ VPWR VGND sg13g2_mux2_1
XFILLER_106_839 VPWR VGND sg13g2_decap_8
XFILLER_105_305 VPWR VGND sg13g2_decap_8
X_06115_ net2961 i_exotiny._0037_\[2\] net1047 _00284_ VPWR VGND sg13g2_mux2_1
X_07095_ net2117 net2289 net914 _00850_ VPWR VGND sg13g2_mux2_1
X_06046_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[18\]
+ net2563 net962 _00231_ VPWR VGND sg13g2_mux2_1
XFILLER_87_712 VPWR VGND sg13g2_fill_1
X_07997_ i_exotiny._2032_ VGND VPWR net532 i_exotiny._2044_\[1\] net1228 sg13g2_dfrbpq_1
XFILLER_86_299 VPWR VGND sg13g2_fill_1
XFILLER_55_620 VPWR VGND sg13g2_fill_2
X_06948_ net2985 net887 _02916_ _02918_ VPWR VGND sg13g2_mux2_1
XFILLER_55_642 VPWR VGND sg13g2_fill_2
X_06879_ net3687 net1094 _02887_ VPWR VGND sg13g2_nor2_1
X_08618_ net1778 VGND VPWR net3673 i_exotiny._1619_\[2\] clknet_leaf_22_clk_regs sg13g2_dfrbpq_2
XFILLER_55_664 VPWR VGND sg13g2_fill_2
XFILLER_54_174 VPWR VGND sg13g2_fill_1
XFILLER_15_539 VPWR VGND sg13g2_fill_1
XFILLER_42_369 VPWR VGND sg13g2_fill_1
X_08549_ net107 VGND VPWR _00623_ i_exotiny._0077_\[0\] clknet_leaf_160_clk_regs sg13g2_dfrbpq_1
X_08618__1358 VPWR VGND net1778 sg13g2_tiehi
XFILLER_24_54 VPWR VGND sg13g2_fill_1
XFILLER_3_900 VPWR VGND sg13g2_decap_8
XFILLER_40_64 VPWR VGND sg13g2_fill_2
XFILLER_2_432 VPWR VGND sg13g2_fill_2
XFILLER_97_509 VPWR VGND sg13g2_decap_8
XFILLER_3_977 VPWR VGND sg13g2_decap_8
X_07936__712 VPWR VGND net712 sg13g2_tiehi
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_18_300 VPWR VGND sg13g2_fill_1
XFILLER_33_325 VPWR VGND sg13g2_fill_2
XFILLER_102_308 VPWR VGND sg13g2_decap_8
X_08256__421 VPWR VGND net421 sg13g2_tiehi
X_07920_ net728 VGND VPWR net1954 i_exotiny._1924_\[13\] clknet_leaf_35_clk_regs sg13g2_dfrbpq_1
XFILLER_68_200 VPWR VGND sg13g2_fill_2
Xhold1906 i_exotiny.i_wb_regs.spi_size_o\[0\] VPWR VGND net3733 sg13g2_dlygate4sd3_1
XFILLER_57_907 VPWR VGND sg13g2_fill_1
Xhold1917 i_exotiny.gpo\[2\] VPWR VGND net3744 sg13g2_dlygate4sd3_1
X_07851_ net2267 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[27\]
+ net983 _01324_ VPWR VGND sg13g2_mux2_1
X_07782_ i_exotiny._0026_\[3\] net874 _03210_ _03215_ VPWR VGND sg13g2_mux2_1
Xhold1939 i_exotiny.i_rstctl.cnt\[4\] VPWR VGND net3766 sg13g2_dlygate4sd3_1
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
X_06802_ _02822_ i_exotiny.i_wb_regs.spi_size_o\[1\] _02745_ VPWR VGND sg13g2_nand2_1
Xhold1928 _00009_ VPWR VGND net3755 sg13g2_dlygate4sd3_1
X_06733_ VGND VPWR _02761_ _02763_ _02764_ net1130 sg13g2_a21oi_1
XFILLER_49_491 VPWR VGND sg13g2_fill_2
X_04994_ _01724_ VPWR _01726_ VGND net1174 _01705_ sg13g2_o21ai_1
XFILLER_24_303 VPWR VGND sg13g2_fill_1
X_06664_ _02703_ _02688_ _02462_ VPWR VGND sg13g2_nand2b_1
X_08263__414 VPWR VGND net414 sg13g2_tiehi
X_05615_ net2050 net1061 _02282_ VPWR VGND sg13g2_nor2_1
X_08403_ net282 VGND VPWR _00477_ i_exotiny._0035_\[2\] clknet_leaf_98_clk_regs sg13g2_dfrbpq_2
X_06595_ i_exotiny._0314_\[11\] net1163 _02653_ VPWR VGND sg13g2_nor2_1
X_08334_ net344 VGND VPWR net2403 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[4\]
+ clknet_leaf_95_clk_regs sg13g2_dfrbpq_1
X_05546_ _02231_ net1275 i_exotiny._0314_\[19\] VPWR VGND sg13g2_nand2b_1
Xclkbuf_leaf_87_clk_regs clknet_5_30__leaf_clk_regs clknet_leaf_87_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08265_ net1175 VGND VPWR net2088 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.genblk7.g_value.r_value[0]
+ clknet_leaf_37_clk_regs sg13g2_dfrbpq_1
X_05477_ VGND VPWR _02178_ i_exotiny._1757_ net1265 sg13g2_or2_1
X_08196_ net481 VGND VPWR _00277_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[27\]
+ clknet_leaf_69_clk_regs sg13g2_dfrbpq_1
X_07216_ net2432 net1090 _02969_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_16_clk_regs clknet_5_6__leaf_clk_regs clknet_leaf_16_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07147_ net2652 net2174 net1011 _00895_ VPWR VGND sg13g2_mux2_1
XFILLER_106_636 VPWR VGND sg13g2_decap_8
XFILLER_105_102 VPWR VGND sg13g2_decap_8
XFILLER_0_903 VPWR VGND sg13g2_decap_8
X_07078_ net3073 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[10\]
+ net916 _00833_ VPWR VGND sg13g2_mux2_1
XFILLER_105_179 VPWR VGND sg13g2_decap_8
Xfanout1019 _02923_ net1019 VPWR VGND sg13g2_buf_8
X_06029_ _02509_ net1262 _02484_ VPWR VGND sg13g2_nand2_2
Xfanout1008 net1009 net1008 VPWR VGND sg13g2_buf_8
XFILLER_102_853 VPWR VGND sg13g2_decap_8
XFILLER_48_907 VPWR VGND sg13g2_fill_2
XFILLER_101_352 VPWR VGND sg13g2_decap_8
XFILLER_19_98 VPWR VGND sg13g2_fill_1
XFILLER_55_450 VPWR VGND sg13g2_fill_1
XFILLER_35_42 VPWR VGND sg13g2_fill_1
XFILLER_42_133 VPWR VGND sg13g2_decap_4
X_08383__295 VPWR VGND net295 sg13g2_tiehi
XFILLER_100_1001 VPWR VGND sg13g2_decap_8
X_08500__180 VPWR VGND net180 sg13g2_tiehi
XFILLER_83_1007 VPWR VGND sg13g2_decap_8
XFILLER_97_317 VPWR VGND sg13g2_decap_8
XFILLER_3_774 VPWR VGND sg13g2_decap_8
XFILLER_32_8 VPWR VGND sg13g2_fill_1
X_08390__288 VPWR VGND net288 sg13g2_tiehi
XFILLER_93_501 VPWR VGND sg13g2_fill_2
XFILLER_65_269 VPWR VGND sg13g2_fill_2
XFILLER_53_409 VPWR VGND sg13g2_fill_2
XFILLER_18_130 VPWR VGND sg13g2_fill_1
XFILLER_92_70 VPWR VGND sg13g2_fill_1
XFILLER_33_144 VPWR VGND sg13g2_fill_1
XFILLER_34_678 VPWR VGND sg13g2_decap_4
X_05400_ i_exotiny._2034_\[4\] _02113_ _02115_ VPWR VGND sg13g2_and2_1
XFILLER_21_306 VPWR VGND sg13g2_fill_1
XFILLER_33_188 VPWR VGND sg13g2_fill_1
X_06380_ _02570_ net2522 net1029 _00506_ VPWR VGND sg13g2_mux2_1
X_05331_ VGND VPWR _01388_ _02054_ _02055_ _01396_ sg13g2_a21oi_1
X_08050_ net644 VGND VPWR net2434 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[19\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
X_05262_ _01987_ VPWR _01988_ VGND _01982_ _01986_ sg13g2_o21ai_1
X_07001_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[5\]
+ net2089 net920 _00768_ VPWR VGND sg13g2_mux2_1
X_08922__1060 VPWR VGND net1480 sg13g2_tiehi
X_05193_ _01921_ i_exotiny._0024_\[1\] _01789_ VPWR VGND sg13g2_nand2_1
X_08952_ net1450 VGND VPWR _01010_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[18\]
+ clknet_leaf_54_clk_regs sg13g2_dfrbpq_1
XFILLER_102_149 VPWR VGND sg13g2_fill_1
X_08883_ net1519 VGND VPWR net1906 i_exotiny.i_wb_spi.dat_rx_r\[13\] clknet_leaf_59_clk_regs
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_134_clk_regs clknet_5_20__leaf_clk_regs clknet_leaf_134_clk_regs VPWR
+ VGND sg13g2_buf_8
X_07903_ net50 VGND VPWR _00004_ i_exotiny._1308_ clknet_leaf_6_clk_regs sg13g2_dfrbpq_1
XFILLER_99_1003 VPWR VGND sg13g2_decap_8
XFILLER_97_884 VPWR VGND sg13g2_decap_8
XFILLER_96_350 VPWR VGND sg13g2_decap_8
Xhold1725 i_exotiny._1902_\[3\] VPWR VGND net3552 sg13g2_dlygate4sd3_1
Xhold1703 i_exotiny.i_wb_spi.dat_rx_r\[31\] VPWR VGND net3530 sg13g2_dlygate4sd3_1
X_07834_ net2142 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[10\]
+ net984 _01307_ VPWR VGND sg13g2_mux2_1
Xhold1714 i_exotiny._1160_\[16\] VPWR VGND net3541 sg13g2_dlygate4sd3_1
Xhold1736 i_exotiny._1617_\[2\] VPWR VGND net3563 sg13g2_dlygate4sd3_1
Xhold1747 i_exotiny.i_wb_spi.dat_rx_r\[2\] VPWR VGND net3574 sg13g2_dlygate4sd3_1
Xhold1758 i_exotiny._1611_\[7\] VPWR VGND net3585 sg13g2_dlygate4sd3_1
Xhold1769 i_exotiny._0369_\[15\] VPWR VGND net3596 sg13g2_dlygate4sd3_1
X_07765_ net2951 net2241 net992 _01250_ VPWR VGND sg13g2_mux2_1
XFILLER_53_910 VPWR VGND sg13g2_fill_1
X_04977_ net1180 _01708_ _01709_ VPWR VGND sg13g2_nor2_1
XFILLER_44_409 VPWR VGND sg13g2_fill_1
XFILLER_64_280 VPWR VGND sg13g2_fill_2
X_06716_ VGND VPWR _02748_ _02749_ _02750_ net1137 sg13g2_a21oi_1
XFILLER_53_932 VPWR VGND sg13g2_fill_1
X_07696_ net2727 _03196_ net999 _01196_ VPWR VGND sg13g2_mux2_1
XFILLER_13_807 VPWR VGND sg13g2_fill_1
X_06647_ net1268 _01461_ _02440_ _02441_ _02688_ VPWR VGND sg13g2_and4_1
X_06578_ net3382 net1155 _02642_ VPWR VGND sg13g2_nor2_1
X_08317_ net361 VGND VPWR _00398_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[19\]
+ clknet_leaf_73_clk_regs sg13g2_dfrbpq_1
X_09297_ net1769 VGND VPWR net2191 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[23\]
+ clknet_leaf_178_clk_regs sg13g2_dfrbpq_1
X_05529_ VGND VPWR net3498 net1276 _02217_ _02216_ sg13g2_a21oi_1
X_08248_ net429 VGND VPWR net2264 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[15\]
+ clknet_leaf_60_clk_regs sg13g2_dfrbpq_1
X_07926__722 VPWR VGND net722 sg13g2_tiehi
XFILLER_21_895 VPWR VGND sg13g2_fill_2
XFILLER_106_433 VPWR VGND sg13g2_decap_8
X_08179_ net498 VGND VPWR _00260_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[10\]
+ clknet_leaf_70_clk_regs sg13g2_dfrbpq_1
X_08742__1246 VPWR VGND net1666 sg13g2_tiehi
XFILLER_0_777 VPWR VGND sg13g2_decap_8
X_07933__715 VPWR VGND net715 sg13g2_tiehi
XFILLER_90_526 VPWR VGND sg13g2_fill_1
XFILLER_28_483 VPWR VGND sg13g2_fill_1
X_08964__1018 VPWR VGND net1438 sg13g2_tiehi
XFILLER_55_280 VPWR VGND sg13g2_fill_1
XFILLER_102_91 VPWR VGND sg13g2_fill_1
X_08246__431 VPWR VGND net431 sg13g2_tiehi
XFILLER_71_795 VPWR VGND sg13g2_fill_1
X_08718__1270 VPWR VGND net1690 sg13g2_tiehi
X_08253__424 VPWR VGND net424 sg13g2_tiehi
X_04900_ _01614_ _01617_ _01632_ VPWR VGND sg13g2_nor2_2
X_05880_ _02466_ _01837_ _02268_ VPWR VGND sg13g2_nand2_1
X_04831_ _01571_ net3640 _01570_ VPWR VGND sg13g2_nand2_1
X_08613__1363 VPWR VGND net1783 sg13g2_tiehi
X_07550_ net3658 _03137_ _03139_ VPWR VGND sg13g2_and2_1
X_04762_ _01513_ net1265 _01510_ VPWR VGND sg13g2_nand2_2
X_06501_ net2703 net888 _02614_ _02616_ VPWR VGND sg13g2_mux2_1
X_09220_ net759 VGND VPWR _01275_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[10\]
+ clknet_leaf_136_clk_regs sg13g2_dfrbpq_1
X_04693_ net1279 _01370_ _01449_ _01451_ VPWR VGND sg13g2_a21o_2
X_07481_ VGND VPWR _01387_ net903 _01070_ _03107_ sg13g2_a21oi_1
X_08820__1168 VPWR VGND net1588 sg13g2_tiehi
X_06432_ net3721 net3697 _02607_ _00521_ VPWR VGND sg13g2_mux2_1
X_06363_ net2764 net2292 net1032 _00493_ VPWR VGND sg13g2_mux2_1
X_08260__417 VPWR VGND net417 sg13g2_tiehi
X_09151_ net831 VGND VPWR net3177 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[7\]
+ clknet_leaf_172_clk_regs sg13g2_dfrbpq_1
X_09082_ net1320 VGND VPWR net2463 i_exotiny._0024_\[2\] clknet_leaf_142_clk_regs
+ sg13g2_dfrbpq_2
X_05314_ net1109 _02038_ _02040_ VPWR VGND sg13g2_nor2_1
X_08102_ net592 VGND VPWR net2441 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[7\]
+ clknet_leaf_126_clk_regs sg13g2_dfrbpq_1
X_08033_ net661 VGND VPWR net2868 i_exotiny._0019_\[2\] clknet_leaf_53_clk_regs sg13g2_dfrbpq_2
X_06294_ net3206 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[26\]
+ net939 _00437_ VPWR VGND sg13g2_mux2_1
Xhold811 _00217_ VPWR VGND net2638 sg13g2_dlygate4sd3_1
X_05245_ _01825_ _01970_ _01971_ _01972_ VPWR VGND sg13g2_nor3_1
Xhold800 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[6\]
+ VPWR VGND net2627 sg13g2_dlygate4sd3_1
X_08438__247 VPWR VGND net247 sg13g2_tiehi
Xhold844 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[30\]
+ VPWR VGND net2671 sg13g2_dlygate4sd3_1
Xhold822 _00536_ VPWR VGND net2649 sg13g2_dlygate4sd3_1
Xhold833 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[29\]
+ VPWR VGND net2660 sg13g2_dlygate4sd3_1
Xhold855 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[29\]
+ VPWR VGND net2682 sg13g2_dlygate4sd3_1
X_05176_ VPWR VGND _01607_ _01901_ _01872_ i_exotiny._0550_ _01904_ _01829_ sg13g2_a221oi_1
XFILLER_104_937 VPWR VGND sg13g2_decap_8
Xhold888 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[16\]
+ VPWR VGND net2715 sg13g2_dlygate4sd3_1
Xhold866 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[24\]
+ VPWR VGND net2693 sg13g2_dlygate4sd3_1
Xhold877 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[30\]
+ VPWR VGND net2704 sg13g2_dlygate4sd3_1
XFILLER_103_458 VPWR VGND sg13g2_decap_8
Xhold899 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[27\]
+ VPWR VGND net2726 sg13g2_dlygate4sd3_1
XFILLER_88_158 VPWR VGND sg13g2_fill_2
Xhold1500 _02106_ VPWR VGND net3327 sg13g2_dlygate4sd3_1
X_08935_ net1467 VGND VPWR _00993_ i_exotiny._0042_\[1\] clknet_leaf_68_clk_regs sg13g2_dfrbpq_2
XFILLER_69_361 VPWR VGND sg13g2_fill_2
XFILLER_69_350 VPWR VGND sg13g2_fill_2
XFILLER_96_180 VPWR VGND sg13g2_fill_2
Xhold1544 _00109_ VPWR VGND net3371 sg13g2_dlygate4sd3_1
X_08866_ net1540 VGND VPWR net2108 i_exotiny.i_wb_regs.spi_cpol_o clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_2
Xhold1522 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[8\]
+ VPWR VGND net3349 sg13g2_dlygate4sd3_1
Xhold1511 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[18\]
+ VPWR VGND net3338 sg13g2_dlygate4sd3_1
Xhold1533 i_exotiny._1160_\[25\] VPWR VGND net3360 sg13g2_dlygate4sd3_1
Xhold1566 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[5\]
+ VPWR VGND net3393 sg13g2_dlygate4sd3_1
Xhold1555 i_exotiny._0314_\[9\] VPWR VGND net3382 sg13g2_dlygate4sd3_1
X_08797_ net1611 VGND VPWR _00855_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[28\]
+ clknet_leaf_167_clk_regs sg13g2_dfrbpq_1
X_07817_ net3375 _03219_ net892 _01294_ VPWR VGND sg13g2_mux2_1
Xhold1577 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[15\]
+ VPWR VGND net3404 sg13g2_dlygate4sd3_1
Xhold1599 _00814_ VPWR VGND net3426 sg13g2_dlygate4sd3_1
X_07748_ net3157 i_exotiny._0026_\[0\] net991 _01233_ VPWR VGND sg13g2_mux2_1
XFILLER_72_537 VPWR VGND sg13g2_decap_4
XFILLER_72_526 VPWR VGND sg13g2_fill_1
Xhold1588 i_exotiny._1160_\[26\] VPWR VGND net3415 sg13g2_dlygate4sd3_1
X_07679_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[14\]
+ net3181 net1001 _01181_ VPWR VGND sg13g2_mux2_1
XFILLER_41_924 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_31_clk_regs clknet_5_8__leaf_clk_regs clknet_leaf_31_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_13_659 VPWR VGND sg13g2_fill_1
XFILLER_12_169 VPWR VGND sg13g2_fill_1
X_08380__298 VPWR VGND net298 sg13g2_tiehi
X_08276__402 VPWR VGND net402 sg13g2_tiehi
XFILLER_10_1012 VPWR VGND sg13g2_decap_8
XFILLER_5_847 VPWR VGND sg13g2_decap_8
XFILLER_106_230 VPWR VGND sg13g2_decap_8
XFILLER_79_103 VPWR VGND sg13g2_fill_1
XFILLER_76_821 VPWR VGND sg13g2_fill_1
XFILLER_57_51 VPWR VGND sg13g2_fill_1
XFILLER_48_545 VPWR VGND sg13g2_fill_1
XFILLER_90_301 VPWR VGND sg13g2_fill_2
XFILLER_29_792 VPWR VGND sg13g2_fill_1
XFILLER_48_589 VPWR VGND sg13g2_fill_2
XFILLER_89_1002 VPWR VGND sg13g2_decap_8
Xhold107 _00937_ VPWR VGND net1934 sg13g2_dlygate4sd3_1
X_09264__101 VPWR VGND net101 sg13g2_tiehi
Xhold118 i_exotiny.i_wb_spi.dat_rx_r\[14\] VPWR VGND net1945 sg13g2_dlygate4sd3_1
X_05030_ _01762_ net1240 VPWR VGND net1238 sg13g2_nand2b_2
Xhold129 _01044_ VPWR VGND net1956 sg13g2_dlygate4sd3_1
XFILLER_99_968 VPWR VGND sg13g2_decap_8
XFILLER_98_467 VPWR VGND sg13g2_decap_8
X_06981_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[23\]
+ net2925 net1019 _00754_ VPWR VGND sg13g2_mux2_1
X_05932_ _02485_ _02484_ VPWR VGND net1262 sg13g2_nand2b_2
X_08720_ net1688 VGND VPWR _00778_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[15\]
+ clknet_leaf_117_clk_regs sg13g2_dfrbpq_1
Xfanout1191 net1192 net1191 VPWR VGND sg13g2_buf_8
X_08651_ net1746 VGND VPWR net2193 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[20\]
+ clknet_leaf_146_clk_regs sg13g2_dfrbpq_1
XFILLER_14_0 VPWR VGND sg13g2_fill_2
X_05863_ VGND VPWR _02448_ _02450_ _02451_ _02429_ sg13g2_a21oi_1
Xfanout1180 _01707_ net1180 VPWR VGND sg13g2_buf_8
XFILLER_96_1028 VPWR VGND sg13g2_fill_1
X_07602_ VGND VPWR i_exotiny.i_wdg_top.clk_div_inst.cnt\[11\] _03170_ _03172_ net1890
+ sg13g2_a21oi_1
X_07916__732 VPWR VGND net732 sg13g2_tiehi
X_04814_ _01556_ VPWR _10679_/A VGND i_exotiny._1793_ net1218 sg13g2_o21ai_1
X_05794_ _02412_ VPWR _00078_ VGND _00022_ _01551_ sg13g2_o21ai_1
X_08582_ net1818 VGND VPWR _00655_ i_exotiny._0314_\[27\] clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
X_04745_ net1254 net1243 _01498_ _01499_ VPWR VGND sg13g2_nor3_2
X_07533_ i_exotiny._1265_ _01474_ net3819 _03128_ VPWR VGND sg13g2_nand3_1
X_04676_ i_exotiny._0327_\[0\] net1234 _01437_ VPWR VGND sg13g2_nor2_2
X_07464_ net1208 _02989_ net3360 _03099_ VPWR VGND sg13g2_nand3_1
X_09203_ net778 VGND VPWR net2697 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[25\]
+ clknet_leaf_79_clk_regs sg13g2_dfrbpq_1
X_06415_ i_exotiny._0327_\[0\] net3688 _02596_ _02597_ VPWR VGND sg13g2_nor3_1
X_09134_ net848 VGND VPWR net2500 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[22\]
+ clknet_leaf_156_clk_regs sg13g2_dfrbpq_1
X_07395_ VGND VPWR i_exotiny._1160_\[11\] net1208 _03048_ _03047_ sg13g2_a21oi_1
X_06346_ net3261 net3419 net1029 _00476_ VPWR VGND sg13g2_mux2_1
X_09065_ net1337 VGND VPWR _01120_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[5\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_1
X_06277_ net2832 net2881 net939 _00420_ VPWR VGND sg13g2_mux2_1
Xhold630 _00167_ VPWR VGND net2457 sg13g2_dlygate4sd3_1
X_08016_ net678 VGND VPWR _00097_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[17\]
+ clknet_leaf_68_clk_regs sg13g2_dfrbpq_1
X_07923__725 VPWR VGND net725 sg13g2_tiehi
X_05228_ VGND VPWR _01956_ i_exotiny._0018_\[1\] net1257 sg13g2_or2_1
Xhold663 _00129_ VPWR VGND net2490 sg13g2_dlygate4sd3_1
Xhold641 _00967_ VPWR VGND net2468 sg13g2_dlygate4sd3_1
Xhold652 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[24\]
+ VPWR VGND net2479 sg13g2_dlygate4sd3_1
XFILLER_2_817 VPWR VGND sg13g2_decap_8
XFILLER_104_734 VPWR VGND sg13g2_decap_8
Xhold696 _00506_ VPWR VGND net2523 sg13g2_dlygate4sd3_1
Xhold674 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[19\]
+ VPWR VGND net2501 sg13g2_dlygate4sd3_1
Xhold685 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[25\]
+ VPWR VGND net2512 sg13g2_dlygate4sd3_1
X_05159_ _01889_ _01653_ i_exotiny._0038_\[2\] _01618_ i_exotiny._0031_\[2\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_103_255 VPWR VGND sg13g2_decap_8
XFILLER_89_489 VPWR VGND sg13g2_fill_1
X_08236__441 VPWR VGND net441 sg13g2_tiehi
X_08918_ net1484 VGND VPWR net2310 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[16\]
+ clknet_leaf_63_clk_regs sg13g2_dfrbpq_1
Xhold1330 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[4\]
+ VPWR VGND net3157 sg13g2_dlygate4sd3_1
XFILLER_100_973 VPWR VGND sg13g2_decap_8
XFILLER_85_651 VPWR VGND sg13g2_fill_2
Xhold1341 i_exotiny._0042_\[2\] VPWR VGND net3168 sg13g2_dlygate4sd3_1
Xhold1352 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[4\]
+ VPWR VGND net3179 sg13g2_dlygate4sd3_1
Xhold1374 i_exotiny.i_wdg_top.clk_div_inst.cnt\[1\] VPWR VGND net3201 sg13g2_dlygate4sd3_1
Xhold1385 i_exotiny._0028_\[3\] VPWR VGND net3212 sg13g2_dlygate4sd3_1
X_08849_ net1557 VGND VPWR _00907_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[16\]
+ clknet_leaf_185_clk_regs sg13g2_dfrbpq_1
Xhold1363 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[13\]
+ VPWR VGND net3190 sg13g2_dlygate4sd3_1
XFILLER_17_217 VPWR VGND sg13g2_fill_1
X_08692__1296 VPWR VGND net1716 sg13g2_tiehi
Xhold1396 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[28\]
+ VPWR VGND net3223 sg13g2_dlygate4sd3_1
XFILLER_27_87 VPWR VGND sg13g2_fill_1
XFILLER_72_378 VPWR VGND sg13g2_fill_1
X_07930__718 VPWR VGND net718 sg13g2_tiehi
X_08881__1101 VPWR VGND net1521 sg13g2_tiehi
XFILLER_40_220 VPWR VGND sg13g2_fill_1
XFILLER_41_754 VPWR VGND sg13g2_fill_2
X_08243__434 VPWR VGND net434 sg13g2_tiehi
XFILLER_13_489 VPWR VGND sg13g2_fill_1
X_10673_ net22 net21 VPWR VGND sg13g2_buf_1
Xclkbuf_5_0__f_clk_regs clknet_4_0_0_clk_regs clknet_5_0__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_4_187 VPWR VGND sg13g2_fill_1
XFILLER_68_629 VPWR VGND sg13g2_fill_1
XFILLER_68_61 VPWR VGND sg13g2_fill_2
XFILLER_68_50 VPWR VGND sg13g2_fill_1
XFILLER_96_949 VPWR VGND sg13g2_decap_8
XFILLER_1_894 VPWR VGND sg13g2_decap_8
X_08250__427 VPWR VGND net427 sg13g2_tiehi
XFILLER_48_375 VPWR VGND sg13g2_fill_1
X_08428__257 VPWR VGND net257 sg13g2_tiehi
XFILLER_56_1001 VPWR VGND sg13g2_fill_1
XFILLER_17_773 VPWR VGND sg13g2_fill_1
XFILLER_72_890 VPWR VGND sg13g2_fill_2
XFILLER_17_784 VPWR VGND sg13g2_fill_2
XFILLER_17_795 VPWR VGND sg13g2_fill_1
X_06200_ net3205 net2629 net947 _00355_ VPWR VGND sg13g2_mux2_1
XFILLER_13_990 VPWR VGND sg13g2_decap_8
XFILLER_31_286 VPWR VGND sg13g2_fill_1
XFILLER_76_2 VPWR VGND sg13g2_fill_1
X_07180_ _02954_ net1285 _02953_ VPWR VGND sg13g2_nand2_1
X_06131_ net2261 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[18\]
+ net1045 _00300_ VPWR VGND sg13g2_mux2_1
X_06062_ i_exotiny._0025_\[1\] net882 _02510_ _02513_ VPWR VGND sg13g2_mux2_1
X_05013_ VGND VPWR _01743_ _01744_ _01745_ _01702_ sg13g2_a21oi_1
XFILLER_98_264 VPWR VGND sg13g2_decap_8
XFILLER_100_214 VPWR VGND sg13g2_fill_2
XFILLER_100_203 VPWR VGND sg13g2_decap_8
X_08703_ net1705 VGND VPWR _00761_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[30\]
+ clknet_leaf_105_clk_regs sg13g2_dfrbpq_1
X_06964_ net2243 net3372 net1022 _00737_ VPWR VGND sg13g2_mux2_1
XFILLER_104_59 VPWR VGND sg13g2_fill_1
XFILLER_100_269 VPWR VGND sg13g2_decap_8
XFILLER_95_982 VPWR VGND sg13g2_decap_8
X_05915_ net2357 net2693 net975 _00132_ VPWR VGND sg13g2_mux2_1
X_06895_ _02899_ net3422 net1068 VPWR VGND sg13g2_nand2_1
XFILLER_27_526 VPWR VGND sg13g2_decap_4
X_08634_ net1763 VGND VPWR _00702_ i_exotiny._0029_\[3\] clknet_leaf_146_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_27_559 VPWR VGND sg13g2_fill_1
X_05846_ VGND VPWR _02051_ _02265_ _02435_ _02428_ sg13g2_a21oi_1
X_05777_ _02402_ i_exotiny._2034_\[6\] net1127 VPWR VGND sg13g2_nand2_1
X_08266__412 VPWR VGND net412 sg13g2_tiehi
X_08565_ net74 VGND VPWR net3463 i_exotiny._0314_\[10\] clknet_leaf_166_clk_regs sg13g2_dfrbpq_1
XFILLER_42_507 VPWR VGND sg13g2_decap_4
XFILLER_23_721 VPWR VGND sg13g2_fill_1
X_07516_ _01499_ _02437_ _03115_ VPWR VGND sg13g2_nor2_1
XFILLER_35_581 VPWR VGND sg13g2_fill_2
X_04728_ i_exotiny._1309_ _01464_ _01484_ VPWR VGND sg13g2_and2_1
X_08496_ net184 VGND VPWR net2449 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[16\]
+ clknet_leaf_108_clk_regs sg13g2_dfrbpq_1
X_08677__1311 VPWR VGND net1731 sg13g2_tiehi
X_07447_ _03087_ VPWR _01056_ VGND net1081 _03086_ sg13g2_o21ai_1
X_04659_ net1252 net1250 _01420_ VPWR VGND sg13g2_nor2b_2
X_07378_ net1989 _02991_ _03034_ VPWR VGND sg13g2_nor2_1
X_06329_ net2719 net2000 net1033 _00466_ VPWR VGND sg13g2_mux2_1
X_09117_ net865 VGND VPWR _01172_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[5\]
+ clknet_leaf_155_clk_regs sg13g2_dfrbpq_1
X_09048_ net804 VGND VPWR net3391 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r[0]
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
Xhold471 i_exotiny.i_rstctl.cnt\[2\] VPWR VGND net2298 sg13g2_dlygate4sd3_1
Xhold460 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[23\]
+ VPWR VGND net2287 sg13g2_dlygate4sd3_1
X_08273__405 VPWR VGND net405 sg13g2_tiehi
Xhold493 _00148_ VPWR VGND net2320 sg13g2_dlygate4sd3_1
Xhold482 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[20\]
+ VPWR VGND net2309 sg13g2_dlygate4sd3_1
XFILLER_104_597 VPWR VGND sg13g2_fill_2
XFILLER_104_586 VPWR VGND sg13g2_decap_8
Xfanout951 net954 net951 VPWR VGND sg13g2_buf_8
Xfanout940 net941 net940 VPWR VGND sg13g2_buf_1
Xfanout973 net976 net973 VPWR VGND sg13g2_buf_8
Xfanout995 net996 net995 VPWR VGND sg13g2_buf_8
Xfanout962 net965 net962 VPWR VGND sg13g2_buf_8
XFILLER_38_42 VPWR VGND sg13g2_fill_1
Xfanout984 net985 net984 VPWR VGND sg13g2_buf_8
Xhold1160 _00387_ VPWR VGND net2987 sg13g2_dlygate4sd3_1
Xhold1193 _00563_ VPWR VGND net3020 sg13g2_dlygate4sd3_1
Xhold1182 i_exotiny._0030_\[3\] VPWR VGND net3009 sg13g2_dlygate4sd3_1
Xhold1171 i_exotiny._1611_\[21\] VPWR VGND net2998 sg13g2_dlygate4sd3_1
X_08997__985 VPWR VGND net1405 sg13g2_tiehi
XFILLER_41_562 VPWR VGND sg13g2_fill_2
XFILLER_70_62 VPWR VGND sg13g2_fill_1
X_08837__1149 VPWR VGND net1569 sg13g2_tiehi
XFILLER_103_1021 VPWR VGND sg13g2_decap_8
Xclkload16 clkload16/Y clknet_leaf_115_clk_regs VPWR VGND sg13g2_inv_8
XFILLER_6_920 VPWR VGND sg13g2_decap_8
Xclkload27 VPWR clkload27/Y clknet_leaf_24_clk_regs VGND sg13g2_inv_1
Xclkload38 VPWR clkload38/Y clknet_leaf_124_clk_regs VGND sg13g2_inv_1
XFILLER_6_997 VPWR VGND sg13g2_decap_8
XFILLER_95_223 VPWR VGND sg13g2_fill_1
XFILLER_83_407 VPWR VGND sg13g2_fill_1
XFILLER_77_960 VPWR VGND sg13g2_fill_1
X_08755__1233 VPWR VGND net1653 sg13g2_tiehi
XFILLER_92_963 VPWR VGND sg13g2_decap_8
X_05700_ net1117 net1920 _02346_ VPWR VGND sg13g2_nor2b_1
X_06680_ _02714_ _02715_ _02716_ _02717_ VPWR VGND sg13g2_nor3_2
X_05631_ net1943 net1065 _02294_ VPWR VGND sg13g2_nor2_1
X_07913__735 VPWR VGND net735 sg13g2_tiehi
X_08350_ net328 VGND VPWR _00431_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[20\]
+ clknet_leaf_95_clk_regs sg13g2_dfrbpq_1
XFILLER_51_315 VPWR VGND sg13g2_fill_2
X_07301_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[26\]
+ net2290 net908 _01018_ VPWR VGND sg13g2_mux2_1
XFILLER_51_359 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_159_clk_regs clknet_5_7__leaf_clk_regs clknet_leaf_159_clk_regs VPWR
+ VGND sg13g2_buf_8
X_05562_ _02241_ VPWR i_exotiny._1611_\[31\] VGND net1076 _02243_ sg13g2_o21ai_1
X_08281_ net397 VGND VPWR net3189 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[15\]
+ clknet_leaf_100_clk_regs sg13g2_dfrbpq_1
XFILLER_60_893 VPWR VGND sg13g2_fill_1
X_05493_ VGND VPWR i_exotiny._0314_\[3\] net1279 _02190_ _02189_ sg13g2_a21oi_1
X_07232_ net3623 net3646 net1092 _00957_ VPWR VGND sg13g2_mux2_1
X_08226__451 VPWR VGND net451 sg13g2_tiehi
XFILLER_20_768 VPWR VGND sg13g2_fill_1
XFILLER_32_595 VPWR VGND sg13g2_fill_1
X_07163_ net2711 net3167 net1012 _00911_ VPWR VGND sg13g2_mux2_1
X_08977__1005 VPWR VGND net1425 sg13g2_tiehi
X_06114_ net2317 i_exotiny._0037_\[1\] net1047 _00283_ VPWR VGND sg13g2_mux2_1
XFILLER_106_818 VPWR VGND sg13g2_decap_8
X_07094_ net3440 net3464 net916 _00849_ VPWR VGND sg13g2_mux2_1
X_07920__728 VPWR VGND net728 sg13g2_tiehi
X_06045_ net2953 net2604 net961 _00230_ VPWR VGND sg13g2_mux2_1
XFILLER_68_960 VPWR VGND sg13g2_fill_2
X_07996_ net137 VGND VPWR i_exotiny._1611_\[31\] i_exotiny._0369_\[7\] clknet_leaf_15_clk_regs
+ sg13g2_dfrbpq_2
X_08233__444 VPWR VGND net444 sg13g2_tiehi
XFILLER_55_610 VPWR VGND sg13g2_fill_1
X_06947_ net2488 net2575 net927 _00726_ VPWR VGND sg13g2_mux2_1
X_08088__606 VPWR VGND net606 sg13g2_tiehi
X_06878_ VGND VPWR net3422 net1131 _02886_ _02885_ sg13g2_a21oi_1
X_08617_ net1779 VGND VPWR _00689_ i_exotiny._1619_\[1\] clknet_leaf_22_clk_regs sg13g2_dfrbpq_2
X_05829_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[25\]
+ net2543 net1057 _00101_ VPWR VGND sg13g2_mux2_1
X_08548_ net108 VGND VPWR _00622_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[4\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_2
X_08479_ net201 VGND VPWR net3347 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[31\]
+ clknet_leaf_158_clk_regs sg13g2_dfrbpq_1
X_08240__437 VPWR VGND net437 sg13g2_tiehi
XFILLER_10_256 VPWR VGND sg13g2_fill_1
X_08833__1155 VPWR VGND net1575 sg13g2_tiehi
XFILLER_3_956 VPWR VGND sg13g2_decap_8
X_08418__267 VPWR VGND net267 sg13g2_tiehi
X_09296__1351 VPWR VGND net1771 sg13g2_tiehi
XFILLER_105_895 VPWR VGND sg13g2_decap_8
XFILLER_104_383 VPWR VGND sg13g2_decap_8
Xhold290 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[23\]
+ VPWR VGND net2117 sg13g2_dlygate4sd3_1
XFILLER_59_993 VPWR VGND sg13g2_fill_2
XFILLER_65_51 VPWR VGND sg13g2_fill_1
XFILLER_65_40 VPWR VGND sg13g2_fill_1
XFILLER_45_186 VPWR VGND sg13g2_fill_1
XFILLER_53_1004 VPWR VGND sg13g2_fill_1
XFILLER_68_212 VPWR VGND sg13g2_fill_1
XFILLER_96_565 VPWR VGND sg13g2_fill_1
Xhold1907 _02819_ VPWR VGND net3734 sg13g2_dlygate4sd3_1
Xhold1918 _02959_ VPWR VGND net3745 sg13g2_dlygate4sd3_1
X_07850_ net2121 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[26\]
+ net984 _01323_ VPWR VGND sg13g2_mux2_1
Xhold1929 i_exotiny.i_wdg_top.clk_div_inst.cnt\[2\] VPWR VGND net3756 sg13g2_dlygate4sd3_1
X_07781_ _03214_ net3321 net988 _01263_ VPWR VGND sg13g2_mux2_1
X_06801_ VGND VPWR net1099 _02820_ _00676_ _02821_ sg13g2_a21oi_1
XFILLER_56_418 VPWR VGND sg13g2_decap_4
X_04993_ _01704_ _01723_ net1201 _01725_ VPWR VGND sg13g2_nand3_1
X_06732_ _02762_ VPWR _02763_ VGND i_exotiny._0369_\[6\] net1192 sg13g2_o21ai_1
Xinput3 ui_in[1] net3 VPWR VGND sg13g2_buf_1
XFILLER_36_120 VPWR VGND sg13g2_decap_4
XFILLER_37_632 VPWR VGND sg13g2_fill_2
XFILLER_52_613 VPWR VGND sg13g2_fill_2
X_06663_ _02702_ i_exotiny._0314_\[2\] _02262_ VPWR VGND sg13g2_xnor2_1
XFILLER_91_292 VPWR VGND sg13g2_fill_1
X_08402_ net283 VGND VPWR _00476_ i_exotiny._0035_\[1\] clknet_leaf_90_clk_regs sg13g2_dfrbpq_2
X_05614_ VGND VPWR net1067 _02281_ _00029_ _02279_ sg13g2_a21oi_1
XFILLER_52_657 VPWR VGND sg13g2_fill_2
X_06594_ net1198 _02651_ _02652_ _00638_ VPWR VGND sg13g2_nor3_1
X_08333_ net345 VGND VPWR _00414_ i_exotiny._0016_\[3\] clknet_leaf_98_clk_regs sg13g2_dfrbpq_2
X_05545_ _02230_ net3596 net1071 VPWR VGND sg13g2_nand2_1
X_08264_ net413 VGND VPWR _00345_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[31\]
+ clknet_leaf_60_clk_regs sg13g2_dfrbpq_1
X_05476_ _01511_ net1265 _01545_ _02177_ VPWR VGND sg13g2_a21o_1
X_08195_ net482 VGND VPWR _00276_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[26\]
+ clknet_leaf_68_clk_regs sg13g2_dfrbpq_1
X_07215_ net1945 net2432 net1090 _00943_ VPWR VGND sg13g2_mux2_1
XFILLER_106_615 VPWR VGND sg13g2_decap_8
X_07146_ net2079 i_exotiny._0036_\[3\] net1012 _00894_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_56_clk_regs clknet_5_14__leaf_clk_regs clknet_leaf_56_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07077_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[5\]
+ net3039 net916 _00832_ VPWR VGND sg13g2_mux2_1
XFILLER_105_158 VPWR VGND sg13g2_decap_8
X_06028_ VGND VPWR net2012 net1104 _00216_ _02508_ sg13g2_a21oi_1
XFILLER_102_832 VPWR VGND sg13g2_decap_8
XFILLER_99_381 VPWR VGND sg13g2_decap_8
X_08270__408 VPWR VGND net408 sg13g2_tiehi
Xfanout1009 net1010 net1009 VPWR VGND sg13g2_buf_8
X_08987__995 VPWR VGND net1415 sg13g2_tiehi
XFILLER_101_331 VPWR VGND sg13g2_decap_8
XFILLER_0_959 VPWR VGND sg13g2_decap_8
X_07979_ net120 VGND VPWR net3602 i_exotiny._0369_\[17\] clknet_leaf_21_clk_regs sg13g2_dfrbpq_2
XFILLER_56_985 VPWR VGND sg13g2_fill_2
XFILLER_28_676 VPWR VGND sg13g2_fill_2
X_08994__988 VPWR VGND net1408 sg13g2_tiehi
XFILLER_51_64 VPWR VGND sg13g2_fill_1
XFILLER_3_753 VPWR VGND sg13g2_decap_8
XFILLER_2_252 VPWR VGND sg13g2_fill_1
XFILLER_105_692 VPWR VGND sg13g2_decap_8
XFILLER_104_180 VPWR VGND sg13g2_decap_8
X_08216__461 VPWR VGND net461 sg13g2_tiehi
XFILLER_65_259 VPWR VGND sg13g2_fill_1
X_09099__883 VPWR VGND net1303 sg13g2_tiehi
XFILLER_18_153 VPWR VGND sg13g2_fill_1
XFILLER_19_698 VPWR VGND sg13g2_fill_2
X_07910__738 VPWR VGND net738 sg13g2_tiehi
X_05330_ _02052_ _02053_ _01912_ _02054_ VPWR VGND sg13g2_nand3_1
X_08223__454 VPWR VGND net454 sg13g2_tiehi
X_05261_ VGND VPWR net1267 i_exotiny._6090_\[0\] _01987_ _01750_ sg13g2_a21oi_1
X_05192_ _01919_ VPWR _01920_ VGND _01914_ _01918_ sg13g2_o21ai_1
X_07000_ net2059 net2765 net922 _00767_ VPWR VGND sg13g2_mux2_1
X_08078__616 VPWR VGND net616 sg13g2_tiehi
X_08951_ net1451 VGND VPWR _01009_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[17\]
+ clknet_leaf_54_clk_regs sg13g2_dfrbpq_1
XFILLER_102_139 VPWR VGND sg13g2_fill_2
XFILLER_102_128 VPWR VGND sg13g2_fill_2
XFILLER_97_863 VPWR VGND sg13g2_decap_8
X_08882_ net1520 VGND VPWR net1898 i_exotiny.i_wb_spi.dat_rx_r\[12\] clknet_leaf_59_clk_regs
+ sg13g2_dfrbpq_1
X_07902_ net48 VGND VPWR _00000_ i_exotiny._1429_ clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
Xhold1726 i_exotiny.i_wdg_top.o_wb_dat\[1\] VPWR VGND net3553 sg13g2_dlygate4sd3_1
Xhold1704 _00959_ VPWR VGND net3531 sg13g2_dlygate4sd3_1
XFILLER_5_1008 VPWR VGND sg13g2_decap_8
X_07833_ net3333 net3124 net986 _01306_ VPWR VGND sg13g2_mux2_1
Xhold1715 _01053_ VPWR VGND net3542 sg13g2_dlygate4sd3_1
Xhold1759 i_exotiny.i_rstctl.cnt\[1\] VPWR VGND net3586 sg13g2_dlygate4sd3_1
XFILLER_84_546 VPWR VGND sg13g2_fill_1
Xhold1737 _00682_ VPWR VGND net3564 sg13g2_dlygate4sd3_1
Xhold1748 _00931_ VPWR VGND net3575 sg13g2_dlygate4sd3_1
X_07764_ net2837 net3170 net992 _01249_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_174_clk_regs clknet_5_4__leaf_clk_regs clknet_leaf_174_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08230__447 VPWR VGND net447 sg13g2_tiehi
X_04976_ VPWR VGND _01433_ _01393_ _01431_ _01428_ _01708_ _01429_ sg13g2_a221oi_1
Xclkbuf_leaf_103_clk_regs clknet_5_29__leaf_clk_regs clknet_leaf_103_clk_regs VPWR
+ VGND sg13g2_buf_8
X_06715_ _02749_ _02747_ net6 net1182 net3528 VPWR VGND sg13g2_a22oi_1
X_07695_ net3319 net882 _03193_ _03196_ VPWR VGND sg13g2_mux2_1
XFILLER_38_985 VPWR VGND sg13g2_fill_2
X_08085__609 VPWR VGND net609 sg13g2_tiehi
X_06646_ _02687_ net2446 net1152 VPWR VGND sg13g2_nand2_1
X_08408__277 VPWR VGND net277 sg13g2_tiehi
X_06577_ i_exotiny._0314_\[5\] net1162 _02641_ VPWR VGND sg13g2_nor2_1
X_08316_ net362 VGND VPWR net2181 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[18\]
+ clknet_leaf_76_clk_regs sg13g2_dfrbpq_1
X_09296_ net1771 VGND VPWR _01351_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[22\]
+ clknet_leaf_171_clk_regs sg13g2_dfrbpq_1
X_05528_ net1277 net3612 _02216_ VPWR VGND sg13g2_nor2b_1
X_08247_ net430 VGND VPWR _00328_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[14\]
+ clknet_leaf_49_clk_regs sg13g2_dfrbpq_1
X_05459_ i_exotiny._1660_ VPWR _02166_ VGND i_exotiny._1619_\[2\] _02138_ sg13g2_o21ai_1
XFILLER_20_384 VPWR VGND sg13g2_fill_1
XFILLER_106_412 VPWR VGND sg13g2_decap_8
X_08178_ net499 VGND VPWR net2149 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[9\]
+ clknet_leaf_111_clk_regs sg13g2_dfrbpq_1
XFILLER_21_67 VPWR VGND sg13g2_fill_2
X_07129_ net1287 net1852 _00879_ VPWR VGND sg13g2_and2_1
XFILLER_106_489 VPWR VGND sg13g2_decap_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_29_952 VPWR VGND sg13g2_fill_1
XFILLER_44_911 VPWR VGND sg13g2_fill_2
X_08972__1010 VPWR VGND net1430 sg13g2_tiehi
XFILLER_30_126 VPWR VGND sg13g2_fill_1
XFILLER_7_344 VPWR VGND sg13g2_fill_2
XFILLER_7_47 VPWR VGND sg13g2_fill_1
XFILLER_98_616 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_1_clk_regs clknet_5_0__leaf_clk_regs clknet_leaf_1_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_93_310 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_fill_2
XFILLER_94_866 VPWR VGND sg13g2_fill_2
X_04830_ _01564_ _01565_ _01569_ _01570_ VPWR VGND sg13g2_nor3_2
XFILLER_93_332 VPWR VGND sg13g2_decap_8
XFILLER_38_259 VPWR VGND sg13g2_fill_2
XFILLER_94_899 VPWR VGND sg13g2_decap_8
X_04761_ net1265 _01510_ _01512_ VPWR VGND sg13g2_and2_1
XFILLER_19_484 VPWR VGND sg13g2_fill_1
X_06500_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[31\]
+ net2363 net1023 _00581_ VPWR VGND sg13g2_mux2_1
X_07480_ net3820 net903 _03107_ VPWR VGND sg13g2_nor2_1
X_04692_ VGND VPWR _01449_ _01450_ net1279 _01370_ sg13g2_a21oi_2
XFILLER_34_476 VPWR VGND sg13g2_fill_1
X_06431_ net3733 net3717 _02607_ _00520_ VPWR VGND sg13g2_mux2_1
X_06362_ net2473 net3439 net1031 _00492_ VPWR VGND sg13g2_mux2_1
X_09150_ net832 VGND VPWR net2725 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[6\]
+ clknet_leaf_148_clk_regs sg13g2_dfrbpq_1
X_06293_ net2424 net3362 net940 _00436_ VPWR VGND sg13g2_mux2_1
X_08101_ net593 VGND VPWR _00182_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[6\]
+ clknet_leaf_124_clk_regs sg13g2_dfrbpq_1
X_09081_ net1321 VGND VPWR net2187 i_exotiny._0024_\[1\] clknet_leaf_154_clk_regs
+ sg13g2_dfrbpq_2
X_05313_ VPWR VGND _02012_ net1110 _01988_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[0\]
+ _02039_ net1107 sg13g2_a221oi_1
X_08032_ net662 VGND VPWR net2129 i_exotiny._0019_\[1\] clknet_leaf_60_clk_regs sg13g2_dfrbpq_2
X_05244_ _01970_ _01971_ net35 VPWR VGND sg13g2_nor2_2
Xhold812 i_exotiny._0018_\[3\] VPWR VGND net2639 sg13g2_dlygate4sd3_1
Xhold801 _00765_ VPWR VGND net2628 sg13g2_dlygate4sd3_1
Xhold845 _00377_ VPWR VGND net2672 sg13g2_dlygate4sd3_1
Xhold834 _00920_ VPWR VGND net2661 sg13g2_dlygate4sd3_1
Xhold823 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[13\]
+ VPWR VGND net2650 sg13g2_dlygate4sd3_1
X_05175_ _01902_ _01903_ net40 VPWR VGND sg13g2_nor2_1
XFILLER_104_916 VPWR VGND sg13g2_decap_8
Xhold889 _01004_ VPWR VGND net2716 sg13g2_dlygate4sd3_1
Xhold856 _00311_ VPWR VGND net2683 sg13g2_dlygate4sd3_1
Xhold878 _01295_ VPWR VGND net2705 sg13g2_dlygate4sd3_1
Xhold867 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[28\]
+ VPWR VGND net2694 sg13g2_dlygate4sd3_1
XFILLER_103_437 VPWR VGND sg13g2_decap_8
X_08934_ net1468 VGND VPWR net2439 i_exotiny._0042_\[0\] clknet_leaf_75_clk_regs sg13g2_dfrbpq_2
Xhold1501 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[28\]
+ VPWR VGND net3328 sg13g2_dlygate4sd3_1
X_08984__998 VPWR VGND net1418 sg13g2_tiehi
Xhold1523 _00254_ VPWR VGND net3350 sg13g2_dlygate4sd3_1
X_08865_ net1541 VGND VPWR _00923_ i_exotiny.i_wb_regs.spi_auto_cs_o clknet_leaf_34_clk_regs
+ sg13g2_dfrbpq_2
Xhold1512 _01149_ VPWR VGND net3339 sg13g2_dlygate4sd3_1
X_08369__309 VPWR VGND net309 sg13g2_tiehi
Xhold1534 _01062_ VPWR VGND net3361 sg13g2_dlygate4sd3_1
Xhold1567 _00315_ VPWR VGND net3394 sg13g2_dlygate4sd3_1
Xhold1545 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[10\]
+ VPWR VGND net3372 sg13g2_dlygate4sd3_1
Xhold1556 _00633_ VPWR VGND net3383 sg13g2_dlygate4sd3_1
X_08796_ net1612 VGND VPWR net2217 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[27\]
+ clknet_leaf_164_clk_regs sg13g2_dfrbpq_1
X_07816_ i_exotiny._0023_\[1\] net884 _03216_ _03219_ VPWR VGND sg13g2_mux2_1
X_07747_ VGND VPWR net1166 _03211_ _03210_ net1139 sg13g2_a21oi_2
Xhold1578 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[19\]
+ VPWR VGND net3405 sg13g2_dlygate4sd3_1
Xhold1589 _01063_ VPWR VGND net3416 sg13g2_dlygate4sd3_1
X_04959_ VPWR VGND _01433_ _01386_ _01431_ _01428_ _01691_ _01429_ sg13g2_a221oi_1
XFILLER_16_56 VPWR VGND sg13g2_fill_2
X_07678_ net3138 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[17\]
+ net998 _01180_ VPWR VGND sg13g2_mux2_1
XFILLER_41_914 VPWR VGND sg13g2_fill_1
X_08768__1220 VPWR VGND net1640 sg13g2_tiehi
X_06629_ net1965 net1155 _02676_ VPWR VGND sg13g2_nor2_1
XFILLER_25_487 VPWR VGND sg13g2_fill_1
XFILLER_41_936 VPWR VGND sg13g2_fill_2
X_07983__124 VPWR VGND net124 sg13g2_tiehi
XFILLER_32_44 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_71_clk_regs clknet_5_30__leaf_clk_regs clknet_leaf_71_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_5_815 VPWR VGND sg13g2_fill_2
X_09279_ net63 VGND VPWR net2366 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[5\]
+ clknet_leaf_178_clk_regs sg13g2_dfrbpq_1
X_08206__471 VPWR VGND net471 sg13g2_tiehi
XFILLER_5_826 VPWR VGND sg13g2_decap_8
XFILLER_106_2 VPWR VGND sg13g2_fill_1
X_09089__893 VPWR VGND net1313 sg13g2_tiehi
XFILLER_106_286 VPWR VGND sg13g2_decap_8
XFILLER_103_993 VPWR VGND sg13g2_decap_8
XFILLER_57_30 VPWR VGND sg13g2_fill_1
XFILLER_91_836 VPWR VGND sg13g2_fill_2
XFILLER_75_376 VPWR VGND sg13g2_fill_2
X_08213__464 VPWR VGND net464 sg13g2_tiehi
XFILLER_35_218 VPWR VGND sg13g2_fill_1
X_08913__1069 VPWR VGND net1489 sg13g2_tiehi
XFILLER_90_368 VPWR VGND sg13g2_fill_2
X_08068__626 VPWR VGND net626 sg13g2_tiehi
X_09096__886 VPWR VGND net1306 sg13g2_tiehi
XFILLER_32_969 VPWR VGND sg13g2_fill_1
X_08398__538 VPWR VGND net538 sg13g2_tiehi
Xhold108 i_exotiny.i_wb_spi.dat_rx_r\[6\] VPWR VGND net1935 sg13g2_dlygate4sd3_1
Xhold119 _00942_ VPWR VGND net1946 sg13g2_dlygate4sd3_1
X_08220__457 VPWR VGND net457 sg13g2_tiehi
XFILLER_99_947 VPWR VGND sg13g2_decap_8
XFILLER_98_446 VPWR VGND sg13g2_decap_8
X_08075__619 VPWR VGND net619 sg13g2_tiehi
XFILLER_3_380 VPWR VGND sg13g2_fill_2
X_06980_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[22\]
+ net2770 net1020 _00753_ VPWR VGND sg13g2_mux2_1
XFILLER_79_682 VPWR VGND sg13g2_fill_2
X_05931_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[1\] _02418_ _02484_
+ VPWR VGND sg13g2_nor2b_2
Xfanout1192 net1193 net1192 VPWR VGND sg13g2_buf_2
Xfanout1170 net1171 net1170 VPWR VGND sg13g2_buf_8
Xfanout1181 net1183 net1181 VPWR VGND sg13g2_buf_2
X_08650_ net1747 VGND VPWR net2316 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[19\]
+ clknet_leaf_145_clk_regs sg13g2_dfrbpq_1
X_08573__58 VPWR VGND net58 sg13g2_tiehi
X_05862_ VGND VPWR _01979_ _02431_ _02450_ _02449_ sg13g2_a21oi_1
X_07601_ net1205 net3579 _01126_ VPWR VGND sg13g2_nor2_1
X_04813_ VGND VPWR net1226 i_exotiny._1793_ _01556_ _01555_ sg13g2_a21oi_1
X_05793_ _02412_ net1875 net1145 VPWR VGND sg13g2_nand2_1
X_08581_ net1820 VGND VPWR _00654_ i_exotiny._0314_\[26\] clknet_leaf_5_clk_regs sg13g2_dfrbpq_1
X_04744_ _01498_ net1245 _01421_ VPWR VGND sg13g2_nand2_2
XFILLER_34_240 VPWR VGND sg13g2_fill_1
X_07532_ _03127_ _01363_ _03126_ VPWR VGND sg13g2_nand2_1
X_07463_ _03097_ _03098_ _03078_ _01061_ VPWR VGND sg13g2_nand3_1
X_04675_ VGND VPWR i_exotiny._0315_\[8\] net1201 _01436_ _01430_ sg13g2_a21oi_1
X_09202_ net779 VGND VPWR _01257_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[24\]
+ clknet_leaf_78_clk_regs sg13g2_dfrbpq_1
X_06414_ net1146 _02593_ _01447_ _02596_ VPWR VGND sg13g2_nand3_1
X_09133_ net849 VGND VPWR _01188_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[21\]
+ clknet_leaf_154_clk_regs sg13g2_dfrbpq_1
X_07394_ _03047_ _03046_ _02992_ _03045_ _02993_ VPWR VGND sg13g2_a22oi_1
X_06345_ net2138 i_exotiny._0035_\[0\] net1029 _00475_ VPWR VGND sg13g2_mux2_1
X_09064_ net1338 VGND VPWR net3629 i_exotiny.i_wdg_top.clk_div_inst.cnt\[4\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
X_06276_ net2708 net2402 net942 _00419_ VPWR VGND sg13g2_mux2_1
X_08015_ net679 VGND VPWR _00096_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[16\]
+ clknet_leaf_62_clk_regs sg13g2_dfrbpq_1
Xhold620 _00656_ VPWR VGND net2447 sg13g2_dlygate4sd3_1
X_05227_ _01952_ _01953_ _01951_ _01955_ VPWR VGND _01954_ sg13g2_nand4_1
XFILLER_104_713 VPWR VGND sg13g2_decap_8
Xhold631 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[25\]
+ VPWR VGND net2458 sg13g2_dlygate4sd3_1
Xhold653 _00371_ VPWR VGND net2480 sg13g2_dlygate4sd3_1
Xhold642 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[20\]
+ VPWR VGND net2469 sg13g2_dlygate4sd3_1
X_05158_ _01888_ _01648_ i_exotiny._0033_\[2\] _01631_ i_exotiny._0027_\[2\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_103_234 VPWR VGND sg13g2_decap_8
XFILLER_89_435 VPWR VGND sg13g2_fill_1
Xhold675 _00095_ VPWR VGND net2502 sg13g2_dlygate4sd3_1
Xhold697 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[5\]
+ VPWR VGND net2524 sg13g2_dlygate4sd3_1
Xhold664 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[31\]
+ VPWR VGND net2491 sg13g2_dlygate4sd3_1
Xhold686 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[7\]
+ VPWR VGND net2513 sg13g2_dlygate4sd3_1
X_05089_ _01819_ VPWR _01820_ VGND net1250 _01818_ sg13g2_o21ai_1
Xhold2010 i_exotiny._0079_\[0\] VPWR VGND net3837 sg13g2_dlygate4sd3_1
X_08917_ net1485 VGND VPWR net3353 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[15\]
+ clknet_leaf_66_clk_regs sg13g2_dfrbpq_1
Xhold1331 _01233_ VPWR VGND net3158 sg13g2_dlygate4sd3_1
XFILLER_100_952 VPWR VGND sg13g2_decap_8
XFILLER_94_39 VPWR VGND sg13g2_fill_2
Xhold1342 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[31\]
+ VPWR VGND net3169 sg13g2_dlygate4sd3_1
Xhold1320 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[29\]
+ VPWR VGND net3147 sg13g2_dlygate4sd3_1
X_08848_ net1558 VGND VPWR _00906_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[15\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
XFILLER_27_11 VPWR VGND sg13g2_decap_4
XFILLER_40_1028 VPWR VGND sg13g2_fill_1
Xhold1386 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[12\]
+ VPWR VGND net3213 sg13g2_dlygate4sd3_1
Xhold1364 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[8\]
+ VPWR VGND net3191 sg13g2_dlygate4sd3_1
Xhold1353 _00411_ VPWR VGND net3180 sg13g2_dlygate4sd3_1
Xhold1375 i_exotiny._0032_\[1\] VPWR VGND net3202 sg13g2_dlygate4sd3_1
Xhold1397 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[8\]
+ VPWR VGND net3224 sg13g2_dlygate4sd3_1
X_08779_ net1629 VGND VPWR net3365 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[10\]
+ clknet_leaf_163_clk_regs sg13g2_dfrbpq_1
XFILLER_53_582 VPWR VGND sg13g2_fill_2
X_08709__1279 VPWR VGND net1699 sg13g2_tiehi
X_10672_ net22 net20 VPWR VGND sg13g2_buf_1
X_09277__67 VPWR VGND net67 sg13g2_tiehi
XFILLER_96_928 VPWR VGND sg13g2_decap_8
XFILLER_95_438 VPWR VGND sg13g2_fill_2
XFILLER_1_873 VPWR VGND sg13g2_decap_8
XFILLER_103_790 VPWR VGND sg13g2_decap_8
XFILLER_48_332 VPWR VGND sg13g2_fill_2
XFILLER_76_696 VPWR VGND sg13g2_fill_1
XFILLER_63_313 VPWR VGND sg13g2_fill_2
XFILLER_36_538 VPWR VGND sg13g2_fill_1
XFILLER_90_187 VPWR VGND sg13g2_fill_2
XFILLER_32_722 VPWR VGND sg13g2_fill_2
XFILLER_44_582 VPWR VGND sg13g2_decap_4
XFILLER_17_1019 VPWR VGND sg13g2_fill_1
X_08359__319 VPWR VGND net319 sg13g2_tiehi
XFILLER_9_995 VPWR VGND sg13g2_decap_8
X_06130_ net3171 net3038 net1047 _00299_ VPWR VGND sg13g2_mux2_1
X_06061_ _02512_ net2588 net964 _00245_ VPWR VGND sg13g2_mux2_1
X_05012_ VGND VPWR _01744_ _01742_ _01729_ sg13g2_or2_1
XFILLER_63_1028 VPWR VGND sg13g2_fill_1
X_06963_ net2677 net2944 net1018 _00736_ VPWR VGND sg13g2_mux2_1
XFILLER_104_27 VPWR VGND sg13g2_fill_2
XFILLER_100_248 VPWR VGND sg13g2_decap_8
XFILLER_95_961 VPWR VGND sg13g2_decap_8
X_05914_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[19\]
+ net2433 net973 _00131_ VPWR VGND sg13g2_mux2_1
X_08702_ net1706 VGND VPWR _00760_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[29\]
+ clknet_leaf_111_clk_regs sg13g2_dfrbpq_1
XFILLER_54_302 VPWR VGND sg13g2_fill_2
X_06894_ VPWR _00692_ _02898_ VGND sg13g2_inv_1
X_08633_ net1764 VGND VPWR net2409 i_exotiny._0029_\[2\] clknet_leaf_146_clk_regs
+ sg13g2_dfrbpq_2
X_05845_ VGND VPWR _02434_ _02265_ _02051_ sg13g2_or2_1
X_05776_ net3796 VPWR _00071_ VGND net1143 _02400_ sg13g2_o21ai_1
XFILLER_81_143 VPWR VGND sg13g2_fill_1
X_08564_ net76 VGND VPWR _00637_ i_exotiny._0314_\[9\] clknet_leaf_180_clk_regs sg13g2_dfrbpq_1
XFILLER_81_198 VPWR VGND sg13g2_fill_1
X_07515_ _03114_ net2099 net901 VPWR VGND sg13g2_nand2_1
X_04727_ net1196 _01483_ _00003_ VPWR VGND sg13g2_nor2_1
X_08495_ net185 VGND VPWR _00569_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[15\]
+ clknet_leaf_107_clk_regs sg13g2_dfrbpq_1
XFILLER_23_755 VPWR VGND sg13g2_fill_2
X_07446_ VGND VPWR net3686 net1080 _03087_ _03077_ sg13g2_a21oi_1
X_07377_ VGND VPWR net1077 _03033_ _01040_ _03031_ sg13g2_a21oi_1
XFILLER_13_68 VPWR VGND sg13g2_fill_1
X_06328_ net2016 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[22\]
+ net1035 _00465_ VPWR VGND sg13g2_mux2_1
X_09116_ net866 VGND VPWR _01171_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[4\]
+ clknet_leaf_157_clk_regs sg13g2_dfrbpq_1
X_09047_ net1571 VGND VPWR _01104_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[2\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_2
X_06259_ _02548_ net2741 net1040 _00407_ VPWR VGND sg13g2_mux2_1
X_08203__474 VPWR VGND net474 sg13g2_tiehi
Xhold472 _03136_ VPWR VGND net2299 sg13g2_dlygate4sd3_1
Xhold461 _00099_ VPWR VGND net2288 sg13g2_dlygate4sd3_1
Xhold450 _00274_ VPWR VGND net2277 sg13g2_dlygate4sd3_1
XFILLER_2_626 VPWR VGND sg13g2_fill_2
XFILLER_2_648 VPWR VGND sg13g2_fill_2
X_08058__636 VPWR VGND net636 sg13g2_tiehi
XFILLER_78_906 VPWR VGND sg13g2_fill_2
Xhold494 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[9\]
+ VPWR VGND net2321 sg13g2_dlygate4sd3_1
Xhold483 _00976_ VPWR VGND net2310 sg13g2_dlygate4sd3_1
X_09086__896 VPWR VGND net1316 sg13g2_tiehi
Xfanout952 net953 net952 VPWR VGND sg13g2_buf_8
XFILLER_78_939 VPWR VGND sg13g2_fill_1
Xfanout941 net944 net941 VPWR VGND sg13g2_buf_8
Xfanout930 net931 net930 VPWR VGND sg13g2_buf_8
Xfanout974 net976 net974 VPWR VGND sg13g2_buf_1
Xfanout963 net964 net963 VPWR VGND sg13g2_buf_8
Xfanout985 net987 net985 VPWR VGND sg13g2_buf_8
XFILLER_92_408 VPWR VGND sg13g2_fill_2
XFILLER_86_983 VPWR VGND sg13g2_decap_8
Xfanout996 net997 net996 VPWR VGND sg13g2_buf_8
Xhold1150 _01195_ VPWR VGND net2977 sg13g2_dlygate4sd3_1
XFILLER_38_87 VPWR VGND sg13g2_decap_8
Xhold1194 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[18\]
+ VPWR VGND net3021 sg13g2_dlygate4sd3_1
Xhold1172 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[23\]
+ VPWR VGND net2999 sg13g2_dlygate4sd3_1
Xhold1183 i_exotiny._1160_\[2\] VPWR VGND net3010 sg13g2_dlygate4sd3_1
Xhold1161 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[13\]
+ VPWR VGND net2988 sg13g2_dlygate4sd3_1
XFILLER_72_143 VPWR VGND sg13g2_fill_2
XFILLER_33_519 VPWR VGND sg13g2_fill_1
X_07989__130 VPWR VGND net130 sg13g2_tiehi
X_08210__467 VPWR VGND net467 sg13g2_tiehi
X_09093__889 VPWR VGND net1309 sg13g2_tiehi
X_08065__629 VPWR VGND net629 sg13g2_tiehi
XFILLER_103_1000 VPWR VGND sg13g2_decap_8
X_08845__1141 VPWR VGND net1561 sg13g2_tiehi
Xclkload17 clkload17/Y clknet_leaf_159_clk_regs VPWR VGND sg13g2_inv_2
Xclkload28 clkload28/Y clknet_leaf_50_clk_regs VPWR VGND sg13g2_inv_2
Xclkload39 VPWR clkload39/Y clknet_leaf_67_clk_regs VGND sg13g2_inv_1
XFILLER_6_976 VPWR VGND sg13g2_decap_8
X_08434__251 VPWR VGND net251 sg13g2_tiehi
XFILLER_95_279 VPWR VGND sg13g2_decap_8
XFILLER_92_942 VPWR VGND sg13g2_decap_8
X_05630_ VGND VPWR net1065 _02292_ _00033_ _02293_ sg13g2_a21oi_1
XFILLER_64_699 VPWR VGND sg13g2_fill_1
X_07300_ net2103 net2880 net908 _01017_ VPWR VGND sg13g2_mux2_1
XFILLER_51_349 VPWR VGND sg13g2_fill_1
X_08650__1327 VPWR VGND net1747 sg13g2_tiehi
X_05561_ VGND VPWR net3155 net1275 _02243_ _02242_ sg13g2_a21oi_1
X_08280_ net398 VGND VPWR _00361_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[14\]
+ clknet_leaf_103_clk_regs sg13g2_dfrbpq_1
X_08441__244 VPWR VGND net244 sg13g2_tiehi
X_08796__1192 VPWR VGND net1612 sg13g2_tiehi
X_05492_ net1274 _01390_ _02189_ VPWR VGND sg13g2_nor2_1
X_07231_ net3616 net3623 net1086 _00956_ VPWR VGND sg13g2_mux2_1
XFILLER_74_0 VPWR VGND sg13g2_fill_1
X_07162_ net2442 net3016 net1008 _00910_ VPWR VGND sg13g2_mux2_1
X_06113_ net3111 i_exotiny._0037_\[0\] net1043 _00282_ VPWR VGND sg13g2_mux2_1
XFILLER_30_1027 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_128_clk_regs clknet_5_21__leaf_clk_regs clknet_leaf_128_clk_regs VPWR
+ VGND sg13g2_buf_8
X_07093_ net2158 net2512 net915 _00848_ VPWR VGND sg13g2_mux2_1
X_06044_ net2220 net2240 net961 _00229_ VPWR VGND sg13g2_mux2_1
XFILLER_101_524 VPWR VGND sg13g2_fill_1
XFILLER_101_513 VPWR VGND sg13g2_decap_8
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
X_07995_ net136 VGND VPWR net3799 i_exotiny._0369_\[6\] clknet_leaf_13_clk_regs sg13g2_dfrbpq_2
Xclkbuf_4_5_0_clk_regs clknet_0_clk_regs clknet_4_5_0_clk_regs VPWR VGND sg13g2_buf_8
X_06946_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[26\]
+ net2927 net925 _00725_ VPWR VGND sg13g2_mux2_1
XFILLER_55_644 VPWR VGND sg13g2_fill_1
XFILLER_55_622 VPWR VGND sg13g2_fill_1
X_06877_ net1128 _02883_ _02884_ _02885_ VPWR VGND sg13g2_nor3_1
X_05828_ net2948 net2453 net1053 _00100_ VPWR VGND sg13g2_mux2_1
X_08616_ net1780 VGND VPWR net3669 i_exotiny._1619_\[0\] clknet_leaf_22_clk_regs sg13g2_dfrbpq_2
XFILLER_55_666 VPWR VGND sg13g2_fill_1
XFILLER_55_699 VPWR VGND sg13g2_decap_4
X_05759_ _02390_ i_exotiny._0315_\[2\] _01465_ VPWR VGND sg13g2_nand2_2
X_08547_ net109 VGND VPWR _00621_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[3\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_2
X_08478_ net202 VGND VPWR _00552_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[30\]
+ clknet_leaf_114_clk_regs sg13g2_dfrbpq_1
X_07429_ i_exotiny._1160_\[19\] net1215 _03074_ VPWR VGND sg13g2_nor2_1
XFILLER_40_22 VPWR VGND sg13g2_decap_4
XFILLER_3_935 VPWR VGND sg13g2_decap_8
Xhold280 _02955_ VPWR VGND net2107 sg13g2_dlygate4sd3_1
XFILLER_2_434 VPWR VGND sg13g2_fill_1
XFILLER_105_874 VPWR VGND sg13g2_decap_8
XFILLER_104_362 VPWR VGND sg13g2_decap_8
Xhold291 _00846_ VPWR VGND net2118 sg13g2_dlygate4sd3_1
XFILLER_1_49 VPWR VGND sg13g2_decap_8
X_08349__329 VPWR VGND net329 sg13g2_tiehi
XFILLER_45_121 VPWR VGND sg13g2_decap_8
XFILLER_27_891 VPWR VGND sg13g2_fill_1
XFILLER_33_327 VPWR VGND sg13g2_fill_1
XFILLER_61_669 VPWR VGND sg13g2_fill_2
XFILLER_60_179 VPWR VGND sg13g2_fill_1
XFILLER_53_1027 VPWR VGND sg13g2_fill_2
XFILLER_6_773 VPWR VGND sg13g2_decap_8
XFILLER_6_784 VPWR VGND sg13g2_fill_2
XFILLER_46_4 VPWR VGND sg13g2_decap_8
Xhold1908 i_exotiny.i_wdg_top.o_wb_dat\[0\] VPWR VGND net3735 sg13g2_dlygate4sd3_1
X_07780_ net3270 net878 _03210_ _03214_ VPWR VGND sg13g2_mux2_1
X_06800_ net2063 net1099 _02821_ VPWR VGND sg13g2_nor2_1
Xhold1919 _00927_ VPWR VGND net3746 sg13g2_dlygate4sd3_1
X_08704__1284 VPWR VGND net1704 sg13g2_tiehi
X_04992_ i_exotiny._6090_\[3\] i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data[0]
+ net1180 _01724_ VPWR VGND sg13g2_mux2_1
Xinput4 ui_in[2] net4 VPWR VGND sg13g2_buf_1
X_06731_ VGND VPWR _01409_ net1192 _02762_ net1169 sg13g2_a21oi_1
XFILLER_37_655 VPWR VGND sg13g2_fill_1
X_08401_ net284 VGND VPWR net2139 i_exotiny._0035_\[0\] clknet_leaf_96_clk_regs sg13g2_dfrbpq_2
XFILLER_64_474 VPWR VGND sg13g2_fill_2
X_06662_ VGND VPWR _02696_ _02701_ _00657_ net1194 sg13g2_a21oi_1
XFILLER_18_880 VPWR VGND sg13g2_fill_1
XFILLER_91_282 VPWR VGND sg13g2_fill_2
X_05613_ VGND VPWR i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data[0]
+ net1119 _02281_ _02280_ sg13g2_a21oi_1
X_06593_ net3462 net1156 _02652_ VPWR VGND sg13g2_nor2_1
X_08332_ net346 VGND VPWR net3027 i_exotiny._0016_\[2\] clknet_leaf_107_clk_regs sg13g2_dfrbpq_2
X_05544_ _02227_ VPWR i_exotiny._1611_\[26\] VGND net1074 _02229_ sg13g2_o21ai_1
X_08263_ net414 VGND VPWR net3162 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[30\]
+ clknet_leaf_49_clk_regs sg13g2_dfrbpq_1
X_08048__646 VPWR VGND net646 sg13g2_tiehi
X_07214_ _02968_ VPWR _00942_ VGND _01415_ net1089 sg13g2_o21ai_1
X_08926__1056 VPWR VGND net1476 sg13g2_tiehi
X_05475_ net1076 VPWR i_exotiny._1611_\[5\] VGND _02175_ _02176_ sg13g2_o21ai_1
X_08194_ net483 VGND VPWR net2401 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[25\]
+ clknet_leaf_112_clk_regs sg13g2_dfrbpq_1
X_07145_ net3281 net3397 net1012 _00893_ VPWR VGND sg13g2_mux2_1
X_07076_ net3000 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[8\]
+ net914 _00831_ VPWR VGND sg13g2_mux2_1
XFILLER_105_137 VPWR VGND sg13g2_decap_8
X_08094__600 VPWR VGND net600 sg13g2_tiehi
X_06027_ _00023_ net1104 _02508_ VPWR VGND sg13g2_nor2_1
X_08200__477 VPWR VGND net477 sg13g2_tiehi
XFILLER_102_811 VPWR VGND sg13g2_decap_8
XFILLER_99_360 VPWR VGND sg13g2_decap_8
XFILLER_0_938 VPWR VGND sg13g2_decap_8
XFILLER_101_310 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_96_clk_regs clknet_5_29__leaf_clk_regs clknet_leaf_96_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_48_909 VPWR VGND sg13g2_fill_1
X_09083__899 VPWR VGND net1319 sg13g2_tiehi
XFILLER_102_888 VPWR VGND sg13g2_decap_8
X_08055__639 VPWR VGND net639 sg13g2_tiehi
Xclkbuf_leaf_25_clk_regs clknet_5_9__leaf_clk_regs clknet_leaf_25_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07978_ net119 VGND VPWR net3585 i_exotiny._1840_\[11\] clknet_leaf_16_clk_regs sg13g2_dfrbpq_2
XFILLER_101_387 VPWR VGND sg13g2_decap_8
X_06929_ net2856 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[13\]
+ net924 _00708_ VPWR VGND sg13g2_mux2_1
XFILLER_83_761 VPWR VGND sg13g2_fill_1
XFILLER_55_441 VPWR VGND sg13g2_decap_8
XFILLER_76_1027 VPWR VGND sg13g2_fill_2
XFILLER_16_839 VPWR VGND sg13g2_fill_2
XFILLER_42_102 VPWR VGND sg13g2_decap_4
XFILLER_24_850 VPWR VGND sg13g2_fill_1
X_08424__261 VPWR VGND net261 sg13g2_tiehi
XFILLER_51_32 VPWR VGND sg13g2_fill_2
XFILLER_13_1011 VPWR VGND sg13g2_decap_8
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_105_671 VPWR VGND sg13g2_decap_8
XFILLER_76_40 VPWR VGND sg13g2_fill_2
X_08431__254 VPWR VGND net254 sg13g2_tiehi
XFILLER_46_485 VPWR VGND sg13g2_fill_1
XFILLER_46_496 VPWR VGND sg13g2_fill_2
X_05260_ _01385_ VPWR _01986_ VGND _01984_ _01985_ sg13g2_o21ai_1
X_05191_ VGND VPWR net1267 i_exotiny._6090_\[1\] _01919_ _01750_ sg13g2_a21oi_1
X_08950_ net1452 VGND VPWR net2246 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[16\]
+ clknet_leaf_75_clk_regs sg13g2_dfrbpq_1
XFILLER_97_842 VPWR VGND sg13g2_decap_8
X_08881_ net1521 VGND VPWR _00939_ i_exotiny.i_wb_spi.dat_rx_r\[11\] clknet_leaf_58_clk_regs
+ sg13g2_dfrbpq_1
X_08617__1359 VPWR VGND net1779 sg13g2_tiehi
X_07901_ net47 VGND VPWR _00003_ i_exotiny._1309_ clknet_leaf_12_clk_regs sg13g2_dfrbpq_2
X_08625__1350 VPWR VGND net1770 sg13g2_tiehi
Xhold1716 _00021_ VPWR VGND net3543 sg13g2_dlygate4sd3_1
XFILLER_57_717 VPWR VGND sg13g2_fill_2
X_07832_ net2808 net3119 net986 _01305_ VPWR VGND sg13g2_mux2_1
Xhold1705 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[5\]
+ VPWR VGND net3532 sg13g2_dlygate4sd3_1
XFILLER_96_385 VPWR VGND sg13g2_decap_8
Xhold1727 _00067_ VPWR VGND net3554 sg13g2_dlygate4sd3_1
Xhold1749 i_exotiny.i_wb_spi.dat_rx_r\[1\] VPWR VGND net3576 sg13g2_dlygate4sd3_1
Xhold1738 i_exotiny._1160_\[18\] VPWR VGND net3565 sg13g2_dlygate4sd3_1
X_07763_ net2780 net2743 net990 _01248_ VPWR VGND sg13g2_mux2_1
X_04975_ VPWR VGND _01433_ _01391_ _01431_ _01428_ _01707_ _01429_ sg13g2_a221oi_1
XFILLER_64_260 VPWR VGND sg13g2_fill_2
X_06714_ _02748_ _02746_ net1173 _02745_ net3430 VPWR VGND sg13g2_a22oi_1
X_07694_ net2976 _03195_ net1000 _01195_ VPWR VGND sg13g2_mux2_1
XFILLER_37_474 VPWR VGND sg13g2_fill_1
XFILLER_64_282 VPWR VGND sg13g2_fill_1
X_06645_ net1198 _02685_ _02686_ _00655_ VPWR VGND sg13g2_nor3_1
X_08315_ net363 VGND VPWR _00396_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[17\]
+ clknet_leaf_83_clk_regs sg13g2_dfrbpq_1
Xclkbuf_leaf_143_clk_regs clknet_5_19__leaf_clk_regs clknet_leaf_143_clk_regs VPWR
+ VGND sg13g2_buf_8
X_06576_ net1194 _02639_ _02640_ _00632_ VPWR VGND sg13g2_nor3_1
X_09295_ net1809 VGND VPWR _01350_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[21\]
+ clknet_leaf_177_clk_regs sg13g2_dfrbpq_1
X_05527_ _02215_ net3641 net1069 VPWR VGND sg13g2_nand2_1
X_08246_ net431 VGND VPWR _00327_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[13\]
+ clknet_leaf_48_clk_regs sg13g2_dfrbpq_1
X_05458_ _02163_ _02164_ _02162_ _02165_ VPWR VGND sg13g2_nand3_1
X_08378__300 VPWR VGND net300 sg13g2_tiehi
XFILLER_21_897 VPWR VGND sg13g2_fill_1
X_08177_ net500 VGND VPWR _00258_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[8\]
+ clknet_leaf_111_clk_regs sg13g2_dfrbpq_1
X_07128_ net1287 net1868 _00878_ VPWR VGND sg13g2_and2_1
X_05389_ net1832 _02108_ i_exotiny._2055_\[1\] VPWR VGND sg13g2_nor2_1
X_08339__339 VPWR VGND net339 sg13g2_tiehi
XFILLER_21_57 VPWR VGND sg13g2_fill_1
XFILLER_106_468 VPWR VGND sg13g2_decap_8
X_07059_ net2806 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[25\]
+ net1015 _00820_ VPWR VGND sg13g2_mux2_1
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_101_184 VPWR VGND sg13g2_decap_8
XFILLER_56_750 VPWR VGND sg13g2_fill_2
X_09198__783 VPWR VGND net783 sg13g2_tiehi
XFILLER_15_179 VPWR VGND sg13g2_fill_1
XFILLER_11_330 VPWR VGND sg13g2_fill_2
XFILLER_87_72 VPWR VGND sg13g2_fill_2
X_08038__656 VPWR VGND net656 sg13g2_tiehi
XFILLER_94_878 VPWR VGND sg13g2_decap_8
X_04760_ VPWR _01511_ _01510_ VGND sg13g2_inv_1
XFILLER_61_252 VPWR VGND sg13g2_fill_2
XFILLER_61_241 VPWR VGND sg13g2_fill_2
X_06430_ net1225 _02130_ _02606_ _02607_ VPWR VGND sg13g2_nor3_2
X_04691_ i_exotiny._0315_\[30\] net1278 _01449_ VPWR VGND sg13g2_nor2_1
XFILLER_35_989 VPWR VGND sg13g2_fill_1
X_08084__610 VPWR VGND net610 sg13g2_tiehi
XFILLER_50_937 VPWR VGND sg13g2_fill_2
X_06361_ net2493 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[16\]
+ net1028 _00491_ VPWR VGND sg13g2_mux2_1
X_08045__649 VPWR VGND net649 sg13g2_tiehi
X_06292_ net2383 net2778 net941 _00435_ VPWR VGND sg13g2_mux2_1
X_09080_ net1322 VGND VPWR net3106 i_exotiny._0024_\[0\] clknet_leaf_141_clk_regs
+ sg13g2_dfrbpq_2
X_05312_ _01612_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[0\].i_hadd.a_i
+ _02037_ _02038_ VPWR VGND sg13g2_a21o_2
X_08100_ net594 VGND VPWR net2587 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[5\]
+ clknet_leaf_125_clk_regs sg13g2_dfrbpq_1
X_08031_ net663 VGND VPWR net2483 i_exotiny._0019_\[0\] clknet_leaf_53_clk_regs sg13g2_dfrbpq_2
X_05243_ net1110 _01969_ _01971_ VPWR VGND sg13g2_and2_1
Xhold802 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[8\]
+ VPWR VGND net2629 sg13g2_dlygate4sd3_1
Xhold835 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[24\]
+ VPWR VGND net2662 sg13g2_dlygate4sd3_1
Xhold813 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[31\]
+ VPWR VGND net2640 sg13g2_dlygate4sd3_1
Xhold846 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[31\]
+ VPWR VGND net2673 sg13g2_dlygate4sd3_1
Xhold824 _00456_ VPWR VGND net2651 sg13g2_dlygate4sd3_1
X_05174_ VPWR VGND _01870_ net1109 _01845_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[2\]
+ _01903_ net1107 sg13g2_a221oi_1
XFILLER_103_416 VPWR VGND sg13g2_decap_8
Xhold857 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[8\]
+ VPWR VGND net2684 sg13g2_dlygate4sd3_1
Xhold879 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[15\]
+ VPWR VGND net2706 sg13g2_dlygate4sd3_1
Xhold868 _00851_ VPWR VGND net2695 sg13g2_dlygate4sd3_1
X_08933_ net1469 VGND VPWR _00991_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[31\]
+ clknet_leaf_66_clk_regs sg13g2_dfrbpq_1
X_08091__603 VPWR VGND net603 sg13g2_tiehi
X_08414__271 VPWR VGND net271 sg13g2_tiehi
Xhold1535 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[25\]
+ VPWR VGND net3362 sg13g2_dlygate4sd3_1
Xhold1524 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[4\]
+ VPWR VGND net3351 sg13g2_dlygate4sd3_1
Xhold1502 _00550_ VPWR VGND net3329 sg13g2_dlygate4sd3_1
X_08864_ net1542 VGND VPWR net3438 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[31\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
Xhold1513 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[13\]
+ VPWR VGND net3340 sg13g2_dlygate4sd3_1
XFILLER_84_333 VPWR VGND sg13g2_fill_1
Xhold1546 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[6\]
+ VPWR VGND net3373 sg13g2_dlygate4sd3_1
X_07815_ net3017 _03218_ net893 _01293_ VPWR VGND sg13g2_mux2_1
X_08795_ net1613 VGND VPWR net3465 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[26\]
+ clknet_leaf_169_clk_regs sg13g2_dfrbpq_1
Xhold1568 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[24\]
+ VPWR VGND net3395 sg13g2_dlygate4sd3_1
Xhold1557 i_exotiny._1160_\[24\] VPWR VGND net3384 sg13g2_dlygate4sd3_1
Xhold1579 _00426_ VPWR VGND net3406 sg13g2_dlygate4sd3_1
X_07746_ _02477_ _02564_ _03210_ VPWR VGND sg13g2_nor2_2
X_04958_ _01420_ _01423_ i_exotiny._0315_\[6\] _01690_ VPWR VGND sg13g2_nand3_1
X_07677_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[12\]
+ net2420 net1002 _01179_ VPWR VGND sg13g2_mux2_1
X_04889_ net1256 _01616_ _01620_ _01621_ VPWR VGND sg13g2_nor3_2
X_06628_ i_exotiny._0314_\[22\] net1161 _02675_ VPWR VGND sg13g2_nor2_1
XFILLER_40_436 VPWR VGND sg13g2_fill_2
X_06559_ net3818 net3737 net1216 _00626_ VPWR VGND sg13g2_mux2_1
X_09278_ net65 VGND VPWR _01333_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[4\]
+ clknet_leaf_174_clk_regs sg13g2_dfrbpq_1
X_08421__264 VPWR VGND net264 sg13g2_tiehi
X_08229_ net448 VGND VPWR net3303 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[28\]
+ clknet_leaf_170_clk_regs sg13g2_dfrbpq_1
XFILLER_106_265 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_40_clk_regs clknet_5_10__leaf_clk_regs clknet_leaf_40_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_103_972 VPWR VGND sg13g2_decap_8
XFILLER_90_303 VPWR VGND sg13g2_fill_1
XFILLER_56_591 VPWR VGND sg13g2_fill_2
XFILLER_56_580 VPWR VGND sg13g2_fill_1
X_08921__1061 VPWR VGND net1481 sg13g2_tiehi
XFILLER_44_753 VPWR VGND sg13g2_fill_1
XFILLER_44_764 VPWR VGND sg13g2_fill_1
Xhold109 _00935_ VPWR VGND net1936 sg13g2_dlygate4sd3_1
XFILLER_99_926 VPWR VGND sg13g2_decap_8
XFILLER_98_425 VPWR VGND sg13g2_decap_8
X_05930_ net2430 _02483_ net973 _00143_ VPWR VGND sg13g2_mux2_1
XFILLER_39_503 VPWR VGND sg13g2_fill_1
Xfanout1182 net1183 net1182 VPWR VGND sg13g2_buf_1
Xfanout1171 net1172 net1171 VPWR VGND sg13g2_buf_8
XFILLER_14_2 VPWR VGND sg13g2_fill_1
Xfanout1160 net1162 net1160 VPWR VGND sg13g2_buf_8
X_05861_ _01498_ _01978_ _02449_ VPWR VGND sg13g2_nor2_1
XFILLER_39_547 VPWR VGND sg13g2_fill_1
XFILLER_96_1019 VPWR VGND sg13g2_decap_8
X_07600_ _03171_ net3578 _03170_ VPWR VGND sg13g2_xnor2_1
Xfanout1193 _01450_ net1193 VPWR VGND sg13g2_buf_8
X_08368__310 VPWR VGND net310 sg13g2_tiehi
X_08580_ net1822 VGND VPWR _00653_ i_exotiny._0314_\[25\] clknet_leaf_4_clk_regs sg13g2_dfrbpq_1
X_04812_ VGND VPWR _01555_ i_exotiny._1757_ i_exotiny._1623_ sg13g2_or2_1
X_05792_ _02411_ VPWR _00077_ VGND _00021_ _01551_ sg13g2_o21ai_1
X_07531_ net1270 net1273 net3694 _03126_ VGND VPWR net1893 sg13g2_nor4_2
X_08329__349 VPWR VGND net349 sg13g2_tiehi
X_04743_ net1245 _01421_ _01497_ VPWR VGND sg13g2_and2_1
X_08741__1247 VPWR VGND net1667 sg13g2_tiehi
XFILLER_23_937 VPWR VGND sg13g2_fill_2
X_04674_ _01433_ _01431_ _01430_ _01435_ VPWR VGND sg13g2_a21o_2
X_07462_ _03098_ net1148 _03035_ VPWR VGND sg13g2_nand2_1
X_09201_ net780 VGND VPWR net2520 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[23\]
+ clknet_leaf_77_clk_regs sg13g2_dfrbpq_1
X_06413_ net1219 net1146 _01437_ _02595_ VPWR VGND _02593_ sg13g2_nand4_1
X_07393_ _03046_ _03002_ i_exotiny._1840_\[11\] _03001_ i_exotiny._0369_\[7\] VPWR
+ VGND sg13g2_a22oi_1
X_06344_ VGND VPWR net1140 _02565_ _02566_ net1167 sg13g2_a21oi_1
X_09132_ net850 VGND VPWR net2527 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[20\]
+ clknet_leaf_152_clk_regs sg13g2_dfrbpq_1
X_08990__992 VPWR VGND net1412 sg13g2_tiehi
X_09063_ net1339 VGND VPWR net1887 i_exotiny.i_wdg_top.clk_div_inst.cnt\[3\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
X_06275_ net2385 net2647 net943 _00418_ VPWR VGND sg13g2_mux2_1
X_09188__793 VPWR VGND net793 sg13g2_tiehi
Xhold621 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[16\]
+ VPWR VGND net2448 sg13g2_dlygate4sd3_1
X_08014_ net680 VGND VPWR net2502 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[15\]
+ clknet_leaf_61_clk_regs sg13g2_dfrbpq_1
X_08375__303 VPWR VGND net303 sg13g2_tiehi
Xhold610 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[22\]
+ VPWR VGND net2437 sg13g2_dlygate4sd3_1
X_05226_ _01954_ _01645_ i_exotiny._0025_\[1\] _01625_ i_exotiny._0030_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold654 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[26\]
+ VPWR VGND net2481 sg13g2_dlygate4sd3_1
Xhold632 _00165_ VPWR VGND net2459 sg13g2_dlygate4sd3_1
Xhold643 _01317_ VPWR VGND net2470 sg13g2_dlygate4sd3_1
X_05157_ _01884_ _01885_ _01875_ _01887_ VPWR VGND _01886_ sg13g2_nand4_1
XFILLER_103_213 VPWR VGND sg13g2_decap_8
X_08963__1019 VPWR VGND net1439 sg13g2_tiehi
Xhold676 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[21\]
+ VPWR VGND net2503 sg13g2_dlygate4sd3_1
Xhold665 _00617_ VPWR VGND net2492 sg13g2_dlygate4sd3_1
Xhold687 _00220_ VPWR VGND net2514 sg13g2_dlygate4sd3_1
XFILLER_104_769 VPWR VGND sg13g2_decap_8
Xhold698 _00700_ VPWR VGND net2525 sg13g2_dlygate4sd3_1
Xhold2000 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[3\] VPWR
+ VGND net3827 sg13g2_dlygate4sd3_1
Xhold2011 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r VPWR VGND net3838
+ sg13g2_dlygate4sd3_1
X_05088_ VGND VPWR _01428_ _01431_ _01819_ _01816_ sg13g2_a21oi_1
X_08916_ net1486 VGND VPWR net2340 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[14\]
+ clknet_leaf_64_clk_regs sg13g2_dfrbpq_1
XFILLER_100_931 VPWR VGND sg13g2_decap_8
Xhold1343 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[16\]
+ VPWR VGND net3170 sg13g2_dlygate4sd3_1
XFILLER_85_653 VPWR VGND sg13g2_fill_1
Xhold1332 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[27\]
+ VPWR VGND net3159 sg13g2_dlygate4sd3_1
X_08847_ net1559 VGND VPWR net3215 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[14\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
Xhold1321 _00472_ VPWR VGND net3148 sg13g2_dlygate4sd3_1
Xhold1310 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[11\]
+ VPWR VGND net3137 sg13g2_dlygate4sd3_1
Xhold1365 _00322_ VPWR VGND net3192 sg13g2_dlygate4sd3_1
Xhold1376 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[5\]
+ VPWR VGND net3203 sg13g2_dlygate4sd3_1
Xhold1354 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[18\]
+ VPWR VGND net3181 sg13g2_dlygate4sd3_1
Xhold1387 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[14\]
+ VPWR VGND net3214 sg13g2_dlygate4sd3_1
Xhold1398 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[24\]
+ VPWR VGND net3225 sg13g2_dlygate4sd3_1
X_08778_ net1630 VGND VPWR net2145 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[9\]
+ clknet_leaf_169_clk_regs sg13g2_dfrbpq_1
XFILLER_38_591 VPWR VGND sg13g2_fill_1
X_09195__786 VPWR VGND net786 sg13g2_tiehi
X_07729_ net2517 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[26\]
+ net995 _01225_ VPWR VGND sg13g2_mux2_1
XFILLER_41_701 VPWR VGND sg13g2_fill_1
X_08717__1271 VPWR VGND net1691 sg13g2_tiehi
XFILLER_41_756 VPWR VGND sg13g2_fill_1
X_10671_ net1246 net18 VPWR VGND sg13g2_buf_1
X_08028__666 VPWR VGND net666 sg13g2_tiehi
X_08612__1364 VPWR VGND net1784 sg13g2_tiehi
XFILLER_4_123 VPWR VGND sg13g2_fill_1
X_08939__1043 VPWR VGND net1463 sg13g2_tiehi
XFILLER_96_907 VPWR VGND sg13g2_decap_8
XFILLER_1_852 VPWR VGND sg13g2_decap_8
XFILLER_89_981 VPWR VGND sg13g2_decap_8
X_08074__620 VPWR VGND net620 sg13g2_tiehi
X_08035__659 VPWR VGND net659 sg13g2_tiehi
XFILLER_75_174 VPWR VGND sg13g2_fill_1
XFILLER_84_84 VPWR VGND sg13g2_fill_2
X_08081__613 VPWR VGND net613 sg13g2_tiehi
XFILLER_83_5 VPWR VGND sg13g2_fill_1
XFILLER_20_929 VPWR VGND sg13g2_fill_1
X_08404__281 VPWR VGND net281 sg13g2_tiehi
XFILLER_9_974 VPWR VGND sg13g2_decap_8
X_06060_ i_exotiny._0025_\[0\] net887 _02510_ _02512_ VPWR VGND sg13g2_mux2_1
X_05011_ _01739_ _01742_ _01371_ _01743_ VPWR VGND sg13g2_nand3_1
XFILLER_98_299 VPWR VGND sg13g2_decap_8
X_08759__1229 VPWR VGND net1649 sg13g2_tiehi
X_06962_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[4\]
+ net3309 net1021 _00735_ VPWR VGND sg13g2_mux2_1
XFILLER_104_17 VPWR VGND sg13g2_fill_2
XFILLER_100_227 VPWR VGND sg13g2_decap_8
XFILLER_95_940 VPWR VGND sg13g2_decap_8
X_05913_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[18\]
+ net2123 net974 _00130_ VPWR VGND sg13g2_mux2_1
X_08701_ net1707 VGND VPWR _00759_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[28\]
+ clknet_leaf_104_clk_regs sg13g2_dfrbpq_1
XFILLER_39_322 VPWR VGND sg13g2_fill_2
X_08411__274 VPWR VGND net274 sg13g2_tiehi
X_08632_ net1765 VGND VPWR net2525 i_exotiny._0029_\[1\] clknet_leaf_147_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_39_355 VPWR VGND sg13g2_fill_2
X_06893_ _02898_ _02719_ _02437_ net1068 net3811 VPWR VGND sg13g2_a22oi_1
X_05844_ _02432_ _02430_ _02429_ _02433_ VPWR VGND sg13g2_a21o_1
X_05775_ _02401_ net1126 _01376_ net1145 net3795 VPWR VGND sg13g2_a22oi_1
X_08563_ net78 VGND VPWR _00636_ i_exotiny._0314_\[8\] clknet_leaf_4_clk_regs sg13g2_dfrbpq_1
XFILLER_82_689 VPWR VGND sg13g2_fill_2
X_08494_ net186 VGND VPWR _00568_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[14\]
+ clknet_leaf_93_clk_regs sg13g2_dfrbpq_1
X_07514_ net2024 net3052 net904 _01097_ VPWR VGND sg13g2_mux2_1
X_04726_ VGND VPWR _01435_ _01478_ _01483_ _01482_ sg13g2_a21oi_1
X_07445_ _03086_ net1149 _03018_ net1209 net3637 VPWR VGND sg13g2_a22oi_1
X_04657_ VPWR _01419_ net4 VGND sg13g2_inv_1
X_07376_ _03033_ _03025_ _03032_ net1208 i_exotiny._1160_\[7\] VPWR VGND sg13g2_a22oi_1
X_06327_ net2730 net2113 net1034 _00464_ VPWR VGND sg13g2_mux2_1
X_09115_ net867 VGND VPWR net2634 i_exotiny._0030_\[3\] clknet_leaf_117_clk_regs sg13g2_dfrbpq_2
X_06258_ net3123 net888 _02546_ _02548_ VPWR VGND sg13g2_mux2_1
X_09046_ net1356 VGND VPWR _01103_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[1\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_2
X_05209_ _01921_ _01935_ _01755_ _01937_ VPWR VGND _01936_ sg13g2_nand4_1
X_06189_ _02539_ net2087 net1263 _00346_ VPWR VGND sg13g2_a21o_1
Xhold451 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[22\]
+ VPWR VGND net2278 sg13g2_dlygate4sd3_1
Xhold440 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[31\]
+ VPWR VGND net2267 sg13g2_dlygate4sd3_1
Xhold462 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[27\]
+ VPWR VGND net2289 sg13g2_dlygate4sd3_1
XFILLER_104_544 VPWR VGND sg13g2_fill_2
Xhold473 _01107_ VPWR VGND net2300 sg13g2_dlygate4sd3_1
Xhold495 _00085_ VPWR VGND net2322 sg13g2_dlygate4sd3_1
Xhold484 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[16\]
+ VPWR VGND net2311 sg13g2_dlygate4sd3_1
XFILLER_89_288 VPWR VGND sg13g2_fill_1
Xfanout942 net944 net942 VPWR VGND sg13g2_buf_8
Xfanout931 _02621_ net931 VPWR VGND sg13g2_buf_8
Xfanout920 net923 net920 VPWR VGND sg13g2_buf_8
Xfanout975 net976 net975 VPWR VGND sg13g2_buf_8
Xfanout953 net954 net953 VPWR VGND sg13g2_buf_8
Xfanout964 net965 net964 VPWR VGND sg13g2_buf_8
Xfanout986 net987 net986 VPWR VGND sg13g2_buf_8
Xfanout997 _03200_ net997 VPWR VGND sg13g2_buf_8
Xhold1140 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[16\]
+ VPWR VGND net2967 sg13g2_dlygate4sd3_1
Xhold1151 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[25\]
+ VPWR VGND net2978 sg13g2_dlygate4sd3_1
XFILLER_85_472 VPWR VGND sg13g2_fill_2
XFILLER_57_174 VPWR VGND sg13g2_fill_2
Xhold1162 _00744_ VPWR VGND net2989 sg13g2_dlygate4sd3_1
XFILLER_18_539 VPWR VGND sg13g2_fill_2
Xhold1184 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[26\]
+ VPWR VGND net3011 sg13g2_dlygate4sd3_1
Xhold1173 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[4\]
+ VPWR VGND net3000 sg13g2_dlygate4sd3_1
Xhold1195 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[12\]
+ VPWR VGND net3022 sg13g2_dlygate4sd3_1
XFILLER_61_818 VPWR VGND sg13g2_fill_1
XFILLER_33_509 VPWR VGND sg13g2_fill_1
XFILLER_60_317 VPWR VGND sg13g2_fill_2
XFILLER_26_583 VPWR VGND sg13g2_fill_2
X_08560__84 VPWR VGND net84 sg13g2_tiehi
X_09293__1393 VPWR VGND net1813 sg13g2_tiehi
Xclkload29 VPWR clkload29/Y clknet_leaf_58_clk_regs VGND sg13g2_inv_1
X_08358__320 VPWR VGND net320 sg13g2_tiehi
XFILLER_10_984 VPWR VGND sg13g2_decap_8
XFILLER_6_955 VPWR VGND sg13g2_decap_8
Xclkload18 clknet_leaf_161_clk_regs clkload18/X VPWR VGND sg13g2_buf_8
XFILLER_86_1018 VPWR VGND sg13g2_decap_8
X_08319__359 VPWR VGND net359 sg13g2_tiehi
XFILLER_68_439 VPWR VGND sg13g2_fill_1
XFILLER_64_667 VPWR VGND sg13g2_fill_1
XFILLER_63_133 VPWR VGND sg13g2_fill_2
X_08365__313 VPWR VGND net313 sg13g2_tiehi
XFILLER_92_998 VPWR VGND sg13g2_decap_8
XFILLER_17_572 VPWR VGND sg13g2_fill_1
X_05560_ net1275 net3185 _02242_ VPWR VGND sg13g2_nor2b_1
X_05491_ _02188_ net3387 net1070 VPWR VGND sg13g2_nand2_1
X_07230_ i_exotiny.i_wb_spi.dat_rx_r\[26\] net3616 net1086 _00955_ VPWR VGND sg13g2_mux2_1
X_07161_ net2052 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[18\]
+ net1010 _00909_ VPWR VGND sg13g2_mux2_1
XFILLER_67_0 VPWR VGND sg13g2_fill_1
XFILLER_8_270 VPWR VGND sg13g2_fill_1
X_06112_ VGND VPWR net1165 _02527_ _02526_ net1138 sg13g2_a21oi_2
X_07092_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[20\]
+ net3413 net913 _00847_ VPWR VGND sg13g2_mux2_1
XFILLER_105_319 VPWR VGND sg13g2_decap_8
X_08691__1297 VPWR VGND net1717 sg13g2_tiehi
X_08372__306 VPWR VGND net306 sg13g2_tiehi
X_06043_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[15\]
+ net2611 net963 _00228_ VPWR VGND sg13g2_mux2_1
XFILLER_99_564 VPWR VGND sg13g2_fill_2
X_09185__796 VPWR VGND net796 sg13g2_tiehi
Xclkbuf_leaf_168_clk_regs clknet_5_4__leaf_clk_regs clknet_leaf_168_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08880__1102 VPWR VGND net1522 sg13g2_tiehi
XFILLER_59_417 VPWR VGND sg13g2_fill_1
X_09304__935 VPWR VGND net1355 sg13g2_tiehi
XFILLER_8_1007 VPWR VGND sg13g2_decap_8
X_07994_ net135 VGND VPWR net2736 i_exotiny._0369_\[5\] clknet_leaf_15_clk_regs sg13g2_dfrbpq_2
X_06945_ net2747 net2897 net924 _00724_ VPWR VGND sg13g2_mux2_1
XFILLER_28_815 VPWR VGND sg13g2_fill_2
XFILLER_82_420 VPWR VGND sg13g2_fill_2
X_08018__676 VPWR VGND net676 sg13g2_tiehi
X_06876_ net1172 VPWR _02884_ VGND net3646 net1186 sg13g2_o21ai_1
XFILLER_94_291 VPWR VGND sg13g2_decap_8
X_05827_ net2287 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[19\]
+ net1054 _00099_ VPWR VGND sg13g2_mux2_1
X_08615_ net1781 VGND VPWR net3621 i_exotiny._1616_\[3\] clknet_leaf_20_clk_regs sg13g2_dfrbpq_2
XFILLER_82_464 VPWR VGND sg13g2_fill_2
X_05758_ _01580_ net1992 _00065_ VPWR VGND sg13g2_nor2_1
X_08546_ net110 VGND VPWR _00620_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[2\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_1
X_09192__789 VPWR VGND net789 sg13g2_tiehi
X_05689_ VGND VPWR i_exotiny._1616_\[2\] net1121 _02338_ _02337_ sg13g2_a21oi_1
X_04709_ _01467_ net1253 _01457_ VPWR VGND sg13g2_nand2_2
X_08477_ net203 VGND VPWR _00551_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[29\]
+ clknet_leaf_159_clk_regs sg13g2_dfrbpq_1
X_08064__630 VPWR VGND net630 sg13g2_tiehi
X_09092__890 VPWR VGND net1310 sg13g2_tiehi
X_07428_ VGND VPWR i_exotiny._0369_\[19\] net1147 _03073_ _03052_ sg13g2_a21oi_1
X_07359_ _03020_ _03004_ _02628_ net1079 net3802 VPWR VGND sg13g2_a22oi_1
X_08025__669 VPWR VGND net669 sg13g2_tiehi
XFILLER_3_914 VPWR VGND sg13g2_decap_8
X_09029_ net1373 VGND VPWR _01087_ i_exotiny._0315_\[17\] clknet_leaf_1_clk_regs sg13g2_dfrbpq_2
XFILLER_105_853 VPWR VGND sg13g2_decap_8
XFILLER_104_341 VPWR VGND sg13g2_decap_8
Xhold270 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[8\]
+ VPWR VGND net2097 sg13g2_dlygate4sd3_1
Xhold292 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[5\]
+ VPWR VGND net2119 sg13g2_dlygate4sd3_1
Xhold281 _00924_ VPWR VGND net2108 sg13g2_dlygate4sd3_1
XFILLER_93_718 VPWR VGND sg13g2_fill_2
X_08071__623 VPWR VGND net623 sg13g2_tiehi
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_105_93 VPWR VGND sg13g2_decap_4
XFILLER_105_82 VPWR VGND sg13g2_decap_8
X_08889__1093 VPWR VGND net1513 sg13g2_tiehi
XFILLER_41_361 VPWR VGND sg13g2_fill_2
X_08401__284 VPWR VGND net284 sg13g2_tiehi
XFILLER_39_4 VPWR VGND sg13g2_fill_2
Xhold1909 _00066_ VPWR VGND net3736 sg13g2_dlygate4sd3_1
X_08676__1312 VPWR VGND net1732 sg13g2_tiehi
X_04991_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data[0]
+ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data[0]
+ net1180 _01723_ VPWR VGND sg13g2_mux2_1
XFILLER_77_770 VPWR VGND sg13g2_fill_2
X_06730_ _02761_ net3751 net1183 VPWR VGND sg13g2_nand2_1
Xinput5 ui_in[3] net5 VPWR VGND sg13g2_buf_2
XFILLER_37_634 VPWR VGND sg13g2_fill_1
X_06661_ _02699_ _02691_ _02700_ _02701_ VPWR VGND sg13g2_a21o_1
X_08400_ net285 VGND VPWR net3431 i_exotiny.i_wb_spi.cnt_presc_r\[6\] clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_1
X_05612_ net1119 net1903 _02280_ VPWR VGND sg13g2_nor2b_1
XFILLER_52_659 VPWR VGND sg13g2_fill_1
X_06592_ i_exotiny._0314_\[10\] net1163 _02651_ VPWR VGND sg13g2_nor2_1
X_08331_ net347 VGND VPWR net2120 i_exotiny._0016_\[1\] clknet_leaf_94_clk_regs sg13g2_dfrbpq_2
X_05543_ VGND VPWR net3402 net1276 _02229_ _02228_ sg13g2_a21oi_1
X_08262_ net415 VGND VPWR net3024 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[29\]
+ clknet_leaf_57_clk_regs sg13g2_dfrbpq_1
X_05474_ _02176_ net1284 net3594 VPWR VGND sg13g2_nand2_1
X_07213_ _02968_ net1945 net1090 VPWR VGND sg13g2_nand2_1
X_08193_ net484 VGND VPWR net2277 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[24\]
+ clknet_leaf_110_clk_regs sg13g2_dfrbpq_1
X_07144_ net2204 i_exotiny._0036_\[1\] net1012 _00892_ VPWR VGND sg13g2_mux2_1
XFILLER_105_116 VPWR VGND sg13g2_decap_8
X_07075_ i_exotiny._0015_\[3\] net2359 net916 _00830_ VPWR VGND sg13g2_mux2_1
X_06026_ VGND VPWR net2063 net1103 _00215_ _02507_ sg13g2_a21oi_1
XFILLER_0_917 VPWR VGND sg13g2_decap_8
XFILLER_102_867 VPWR VGND sg13g2_decap_8
XFILLER_101_366 VPWR VGND sg13g2_decap_8
XFILLER_75_707 VPWR VGND sg13g2_decap_8
X_07977_ net118 VGND VPWR i_exotiny._1611_\[6\] i_exotiny._0369_\[30\] clknet_leaf_17_clk_regs
+ sg13g2_dfrbpq_2
X_06928_ net2688 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[12\]
+ net926 _00707_ VPWR VGND sg13g2_mux2_1
X_08348__330 VPWR VGND net330 sg13g2_tiehi
Xclkbuf_leaf_65_clk_regs clknet_5_24__leaf_clk_regs clknet_leaf_65_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06859_ net1129 _02868_ _02869_ _02870_ VPWR VGND sg13g2_nor3_1
XFILLER_56_987 VPWR VGND sg13g2_fill_1
XFILLER_28_678 VPWR VGND sg13g2_fill_1
XFILLER_27_199 VPWR VGND sg13g2_fill_2
X_08529_ net151 VGND VPWR net3055 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[17\]
+ clknet_leaf_176_clk_regs sg13g2_dfrbpq_1
X_08309__369 VPWR VGND net369 sg13g2_tiehi
XFILLER_11_578 VPWR VGND sg13g2_fill_1
XFILLER_100_1015 VPWR VGND sg13g2_decap_8
X_08754__1234 VPWR VGND net1654 sg13g2_tiehi
X_08355__323 VPWR VGND net323 sg13g2_tiehi
XFILLER_105_650 VPWR VGND sg13g2_decap_8
XFILLER_3_788 VPWR VGND sg13g2_decap_8
XFILLER_18_100 VPWR VGND sg13g2_fill_1
X_08976__1006 VPWR VGND net1426 sg13g2_tiehi
XFILLER_18_177 VPWR VGND sg13g2_fill_2
X_08362__316 VPWR VGND net316 sg13g2_tiehi
XFILLER_42_670 VPWR VGND sg13g2_fill_1
X_05190_ _01385_ VPWR _01918_ VGND _01916_ _01917_ sg13g2_o21ai_1
X_09182__799 VPWR VGND net799 sg13g2_tiehi
X_08880_ net1522 VGND VPWR _00938_ i_exotiny.i_wb_spi.dat_rx_r\[10\] clknet_leaf_59_clk_regs
+ sg13g2_dfrbpq_1
X_07900_ net46 VGND VPWR _00002_ i_exotiny._1306_ clknet_leaf_6_clk_regs sg13g2_dfrbpq_2
XFILLER_96_364 VPWR VGND sg13g2_decap_8
Xhold1717 _00214_ VPWR VGND net3544 sg13g2_dlygate4sd3_1
Xhold1706 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[28\]
+ VPWR VGND net3533 sg13g2_dlygate4sd3_1
X_07831_ net3137 net2307 net983 _01304_ VPWR VGND sg13g2_mux2_1
XFILLER_99_1028 VPWR VGND sg13g2_fill_1
XFILLER_99_1017 VPWR VGND sg13g2_decap_8
XFILLER_97_898 VPWR VGND sg13g2_decap_8
X_08054__640 VPWR VGND net640 sg13g2_tiehi
XFILLER_56_228 VPWR VGND sg13g2_fill_2
Xhold1728 i_exotiny._0315_\[9\] VPWR VGND net3555 sg13g2_dlygate4sd3_1
Xhold1739 _01055_ VPWR VGND net3566 sg13g2_dlygate4sd3_1
XFILLER_38_910 VPWR VGND sg13g2_fill_1
X_07762_ net2581 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[14\]
+ net988 _01247_ VPWR VGND sg13g2_mux2_1
X_04974_ net1174 _01705_ _01706_ VPWR VGND sg13g2_nor2_2
X_06713_ _02721_ _02723_ _02747_ VPWR VGND sg13g2_nor2b_2
X_07693_ i_exotiny._0030_\[0\] net887 _03193_ _03195_ VPWR VGND sg13g2_mux2_1
XFILLER_38_987 VPWR VGND sg13g2_fill_1
X_08832__1156 VPWR VGND net1576 sg13g2_tiehi
X_08015__679 VPWR VGND net679 sg13g2_tiehi
X_06644_ net2037 net1154 _02686_ VPWR VGND sg13g2_nor2_1
X_06575_ net3476 net1152 _02640_ VPWR VGND sg13g2_nor2_1
X_08314_ net364 VGND VPWR net2622 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[16\]
+ clknet_leaf_82_clk_regs sg13g2_dfrbpq_1
X_05526_ _02212_ VPWR i_exotiny._1611_\[22\] VGND net1075 _02214_ sg13g2_o21ai_1
X_09294_ net1811 VGND VPWR _01349_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[20\]
+ clknet_leaf_175_clk_regs sg13g2_dfrbpq_1
X_08245_ net432 VGND VPWR net3246 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[12\]
+ clknet_leaf_56_clk_regs sg13g2_dfrbpq_1
X_05457_ _02164_ _02149_ i_exotiny._1617_\[2\] _02148_ i_exotiny._1612_\[2\] VPWR
+ VGND sg13g2_a22oi_1
X_08061__633 VPWR VGND net633 sg13g2_tiehi
X_05388_ VGND VPWR net1112 _02098_ _02108_ _02107_ sg13g2_a21oi_1
X_08176_ net501 VGND VPWR _00257_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[7\]
+ clknet_leaf_69_clk_regs sg13g2_dfrbpq_1
Xclkbuf_leaf_183_clk_regs clknet_5_1__leaf_clk_regs clknet_leaf_183_clk_regs VPWR
+ VGND sg13g2_buf_8
X_07127_ net1287 net1865 _00877_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_112_clk_regs clknet_5_25__leaf_clk_regs clknet_leaf_112_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_21_69 VPWR VGND sg13g2_fill_1
XFILLER_106_447 VPWR VGND sg13g2_decap_8
X_07058_ net3304 net2830 net1013 _00819_ VPWR VGND sg13g2_mux2_1
XFILLER_0_714 VPWR VGND sg13g2_decap_8
XFILLER_88_843 VPWR VGND sg13g2_fill_1
X_06009_ net2630 _02498_ net1049 _00207_ VPWR VGND sg13g2_mux2_1
XFILLER_48_707 VPWR VGND sg13g2_decap_4
XFILLER_87_386 VPWR VGND sg13g2_fill_2
XFILLER_28_442 VPWR VGND sg13g2_fill_1
XFILLER_55_261 VPWR VGND sg13g2_fill_2
XFILLER_44_913 VPWR VGND sg13g2_fill_1
X_08808__1180 VPWR VGND net1600 sg13g2_tiehi
XFILLER_71_754 VPWR VGND sg13g2_fill_2
XFILLER_12_821 VPWR VGND sg13g2_fill_1
XFILLER_30_117 VPWR VGND sg13g2_fill_2
X_08498__182 VPWR VGND net182 sg13g2_tiehi
XFILLER_105_480 VPWR VGND sg13g2_decap_8
XFILLER_94_868 VPWR VGND sg13g2_fill_1
XFILLER_38_239 VPWR VGND sg13g2_fill_2
X_04690_ _01448_ net1270 _01447_ VPWR VGND sg13g2_nand2_1
XFILLER_35_946 VPWR VGND sg13g2_fill_1
XFILLER_50_949 VPWR VGND sg13g2_fill_2
X_06360_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[19\]
+ net2851 net1030 _00490_ VPWR VGND sg13g2_mux2_1
X_06291_ net2887 net2820 net943 _00434_ VPWR VGND sg13g2_mux2_1
X_05311_ _01612_ _02035_ _02036_ _02037_ VPWR VGND sg13g2_nor3_1
X_08030_ net664 VGND VPWR _00111_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[31\]
+ clknet_leaf_62_clk_regs sg13g2_dfrbpq_1
X_05242_ VPWR VGND _01944_ _01607_ _01920_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[1\]
+ _01970_ net1107 sg13g2_a221oi_1
Xhold803 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[31\]
+ VPWR VGND net2630 sg13g2_dlygate4sd3_1
Xhold836 _01016_ VPWR VGND net2663 sg13g2_dlygate4sd3_1
Xhold814 _00410_ VPWR VGND net2641 sg13g2_dlygate4sd3_1
Xhold825 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[8\]
+ VPWR VGND net2652 sg13g2_dlygate4sd3_1
X_05173_ net1109 _01897_ _01902_ VPWR VGND sg13g2_and2_1
Xhold869 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[25\]
+ VPWR VGND net2696 sg13g2_dlygate4sd3_1
X_08338__340 VPWR VGND net340 sg13g2_tiehi
Xhold847 _00438_ VPWR VGND net2674 sg13g2_dlygate4sd3_1
XFILLER_66_1027 VPWR VGND sg13g2_fill_2
Xhold858 _01337_ VPWR VGND net2685 sg13g2_dlygate4sd3_1
X_08932_ net1470 VGND VPWR net2615 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[30\]
+ clknet_leaf_64_clk_regs sg13g2_dfrbpq_1
XFILLER_97_684 VPWR VGND sg13g2_fill_1
Xhold1525 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[15\]
+ VPWR VGND net3352 sg13g2_dlygate4sd3_1
Xhold1514 i_exotiny._0040_\[0\] VPWR VGND net3341 sg13g2_dlygate4sd3_1
X_08863_ net1543 VGND VPWR _00921_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[30\]
+ clknet_leaf_184_clk_regs sg13g2_dfrbpq_1
Xhold1503 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[19\]
+ VPWR VGND net3330 sg13g2_dlygate4sd3_1
Xhold1536 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[12\]
+ VPWR VGND net3363 sg13g2_dlygate4sd3_1
Xhold1547 _00481_ VPWR VGND net3374 sg13g2_dlygate4sd3_1
XFILLER_57_548 VPWR VGND sg13g2_decap_4
X_08794_ net1614 VGND VPWR _00852_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[25\]
+ clknet_leaf_168_clk_regs sg13g2_dfrbpq_1
X_07814_ i_exotiny._0023_\[0\] net887 _03216_ _03218_ VPWR VGND sg13g2_mux2_1
Xhold1558 _01061_ VPWR VGND net3385 sg13g2_dlygate4sd3_1
X_07745_ _03209_ VPWR _01232_ VGND _01397_ net1060 sg13g2_o21ai_1
Xhold1569 _00783_ VPWR VGND net3396 sg13g2_dlygate4sd3_1
X_04957_ _01689_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[1\] _01688_ VPWR
+ VGND sg13g2_nand2_1
XFILLER_25_401 VPWR VGND sg13g2_fill_2
X_07941__85 VPWR VGND net85 sg13g2_tiehi
X_07676_ net2882 net2960 net1001 _01178_ VPWR VGND sg13g2_mux2_1
X_04888_ _01620_ net1260 VPWR VGND net1259 sg13g2_nand2b_2
X_08345__333 VPWR VGND net333 sg13g2_tiehi
X_06627_ net1194 _02673_ _02674_ _00649_ VPWR VGND sg13g2_nor3_1
X_06558_ net3810 net3675 net1216 _00625_ VPWR VGND sg13g2_mux2_1
X_06489_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[20\]
+ net2448 net1026 _00570_ VPWR VGND sg13g2_mux2_1
X_09277_ net67 VGND VPWR _01332_ i_exotiny._0021_\[3\] clknet_leaf_170_clk_regs sg13g2_dfrbpq_2
XFILLER_21_662 VPWR VGND sg13g2_fill_2
X_05509_ VGND VPWR i_exotiny._0314_\[9\] net1275 _02202_ _02201_ sg13g2_a21oi_1
X_08228_ net449 VGND VPWR _00309_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[27\]
+ clknet_leaf_150_clk_regs sg13g2_dfrbpq_1
XFILLER_10_1026 VPWR VGND sg13g2_fill_2
X_08159_ net519 VGND VPWR _00240_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[23\]
+ clknet_leaf_118_clk_regs sg13g2_dfrbpq_1
XFILLER_106_244 VPWR VGND sg13g2_decap_8
XFILLER_103_951 VPWR VGND sg13g2_decap_8
X_08352__326 VPWR VGND net326 sg13g2_tiehi
Xclkbuf_leaf_80_clk_regs clknet_5_27__leaf_clk_regs clknet_leaf_80_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_48_526 VPWR VGND sg13g2_fill_1
XFILLER_102_483 VPWR VGND sg13g2_decap_8
XFILLER_91_838 VPWR VGND sg13g2_fill_1
XFILLER_75_378 VPWR VGND sg13g2_fill_1
XFILLER_106_1021 VPWR VGND sg13g2_decap_8
XFILLER_89_1027 VPWR VGND sg13g2_fill_2
XFILLER_89_1016 VPWR VGND sg13g2_decap_8
X_08044__650 VPWR VGND net650 sg13g2_tiehi
XFILLER_8_666 VPWR VGND sg13g2_fill_2
XFILLER_22_90 VPWR VGND sg13g2_fill_1
XFILLER_99_905 VPWR VGND sg13g2_decap_8
XFILLER_98_404 VPWR VGND sg13g2_decap_8
XFILLER_4_883 VPWR VGND sg13g2_decap_8
XFILLER_100_409 VPWR VGND sg13g2_decap_8
XFILLER_94_621 VPWR VGND sg13g2_fill_2
XFILLER_79_684 VPWR VGND sg13g2_fill_1
Xfanout1150 net1151 net1150 VPWR VGND sg13g2_buf_8
Xfanout1172 net1173 net1172 VPWR VGND sg13g2_buf_1
Xfanout1183 _01515_ net1183 VPWR VGND sg13g2_buf_8
Xfanout1161 net1162 net1161 VPWR VGND sg13g2_buf_1
X_05860_ _01978_ _01979_ _01496_ _02448_ VPWR VGND sg13g2_nand3_1
X_05791_ _02411_ net1870 net1145 VPWR VGND sg13g2_nand2_1
Xfanout1194 net1195 net1194 VPWR VGND sg13g2_buf_8
X_04811_ net1226 _01554_ _00008_ VPWR VGND sg13g2_nor2_1
X_08051__643 VPWR VGND net643 sg13g2_tiehi
X_07530_ _03122_ VPWR _01101_ VGND _03123_ _03125_ sg13g2_o21ai_1
X_04742_ net1243 _01422_ _01496_ VPWR VGND sg13g2_nor2_2
XFILLER_50_702 VPWR VGND sg13g2_fill_2
X_07461_ net1208 _02989_ net3384 _03097_ VPWR VGND sg13g2_nand3_1
X_04673_ _01434_ _01431_ _01433_ _01429_ _01428_ VPWR VGND sg13g2_a22oi_1
XFILLER_97_0 VPWR VGND sg13g2_fill_2
X_09200_ net781 VGND VPWR net2133 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[22\]
+ clknet_leaf_79_clk_regs sg13g2_dfrbpq_1
X_06412_ net1219 net1146 _01437_ _02594_ VPWR VGND sg13g2_nand3_1
X_07392_ _03045_ i_exotiny._0369_\[20\] net1214 VPWR VGND sg13g2_nand2_1
X_06343_ _02532_ _02564_ _02565_ VPWR VGND sg13g2_nor2_2
X_09131_ net851 VGND VPWR net2177 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[19\]
+ clknet_leaf_155_clk_regs sg13g2_dfrbpq_1
X_09062_ net1340 VGND VPWR _01117_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[2\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
X_06274_ net3348 net3026 net939 _00417_ VPWR VGND sg13g2_mux2_1
Xhold611 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[4\]
+ VPWR VGND net2438 sg13g2_dlygate4sd3_1
X_08013_ net681 VGND VPWR net2248 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[14\]
+ clknet_leaf_67_clk_regs sg13g2_dfrbpq_1
Xhold600 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[10\]
+ VPWR VGND net2427 sg13g2_dlygate4sd3_1
X_05225_ _01953_ _01631_ i_exotiny._0027_\[1\] _01626_ i_exotiny._0014_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold633 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[7\]
+ VPWR VGND net2460 sg13g2_dlygate4sd3_1
Xhold622 _00570_ VPWR VGND net2449 sg13g2_dlygate4sd3_1
Xhold644 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[28\]
+ VPWR VGND net2471 sg13g2_dlygate4sd3_1
X_05156_ _01886_ _01655_ i_exotiny._0026_\[2\] _01615_ i_exotiny._0021_\[2\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_104_748 VPWR VGND sg13g2_decap_8
Xhold666 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[20\]
+ VPWR VGND net2493 sg13g2_dlygate4sd3_1
Xhold655 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[4\]
+ VPWR VGND net2482 sg13g2_dlygate4sd3_1
Xhold688 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[23\]
+ VPWR VGND net2515 sg13g2_dlygate4sd3_1
Xhold677 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[22\]
+ VPWR VGND net2504 sg13g2_dlygate4sd3_1
X_08971__1011 VPWR VGND net1431 sg13g2_tiehi
Xhold2012 i_exotiny.i_wdg_top.clk_div_inst.cnt\[19\] VPWR VGND net3839 sg13g2_dlygate4sd3_1
Xhold699 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[24\]
+ VPWR VGND net2526 sg13g2_dlygate4sd3_1
X_05087_ _01818_ net1224 VPWR VGND _01603_ sg13g2_nand2b_2
Xhold2001 i_exotiny._0369_\[20\] VPWR VGND net3828 sg13g2_dlygate4sd3_1
XFILLER_103_269 VPWR VGND sg13g2_decap_8
XFILLER_100_910 VPWR VGND sg13g2_decap_8
XFILLER_98_993 VPWR VGND sg13g2_decap_8
Xhold1300 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[4\]
+ VPWR VGND net3127 sg13g2_dlygate4sd3_1
X_08915_ net1487 VGND VPWR _00973_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[13\]
+ clknet_leaf_113_clk_regs sg13g2_dfrbpq_1
Xhold1322 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[14\]
+ VPWR VGND net3149 sg13g2_dlygate4sd3_1
Xhold1333 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[25\]
+ VPWR VGND net3160 sg13g2_dlygate4sd3_1
X_08846_ net1560 VGND VPWR net2199 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[13\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
Xhold1311 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[13\]
+ VPWR VGND net3138 sg13g2_dlygate4sd3_1
XFILLER_100_987 VPWR VGND sg13g2_decap_8
Xhold1366 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[9\]
+ VPWR VGND net3193 sg13g2_dlygate4sd3_1
Xhold1377 _01266_ VPWR VGND net3204 sg13g2_dlygate4sd3_1
Xhold1344 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[21\]
+ VPWR VGND net3171 sg13g2_dlygate4sd3_1
Xhold1355 _01181_ VPWR VGND net3182 sg13g2_dlygate4sd3_1
X_08488__192 VPWR VGND net192 sg13g2_tiehi
Xhold1388 _00905_ VPWR VGND net3215 sg13g2_dlygate4sd3_1
X_08572__60 VPWR VGND net60 sg13g2_tiehi
Xhold1399 _01285_ VPWR VGND net3226 sg13g2_dlygate4sd3_1
X_08777_ net1631 VGND VPWR _00835_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[8\]
+ clknet_leaf_168_clk_regs sg13g2_dfrbpq_1
X_05989_ net2486 net2395 net1051 _00191_ VPWR VGND sg13g2_mux2_1
XFILLER_45_529 VPWR VGND sg13g2_decap_4
XFILLER_53_551 VPWR VGND sg13g2_decap_4
X_07728_ net2379 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[25\]
+ net997 _01224_ VPWR VGND sg13g2_mux2_1
X_07659_ i_exotiny._0024_\[2\] net879 _03187_ _03191_ VPWR VGND sg13g2_mux2_1
XFILLER_13_426 VPWR VGND sg13g2_fill_1
XFILLER_43_56 VPWR VGND sg13g2_fill_2
X_08495__185 VPWR VGND net185 sg13g2_tiehi
XFILLER_4_28 VPWR VGND sg13g2_decap_4
XFILLER_89_960 VPWR VGND sg13g2_decap_8
XFILLER_1_831 VPWR VGND sg13g2_decap_8
XFILLER_102_280 VPWR VGND sg13g2_decap_8
XFILLER_63_315 VPWR VGND sg13g2_fill_1
XFILLER_1_1013 VPWR VGND sg13g2_decap_8
XFILLER_44_551 VPWR VGND sg13g2_decap_4
X_08328__350 VPWR VGND net350 sg13g2_tiehi
X_08849__1137 VPWR VGND net1557 sg13g2_tiehi
XFILLER_9_920 VPWR VGND sg13g2_fill_1
XFILLER_9_953 VPWR VGND sg13g2_decap_8
X_05010_ _01742_ _01424_ _01741_ VPWR VGND sg13g2_xnor2_1
X_08335__343 VPWR VGND net343 sg13g2_tiehi
XFILLER_98_278 VPWR VGND sg13g2_decap_8
X_08767__1221 VPWR VGND net1641 sg13g2_tiehi
X_06961_ net2805 net3247 net1019 _00734_ VPWR VGND sg13g2_mux2_1
X_05912_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[17\]
+ net2489 net972 _00129_ VPWR VGND sg13g2_mux2_1
X_08700_ net1708 VGND VPWR net2179 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[27\]
+ clknet_leaf_104_clk_regs sg13g2_dfrbpq_1
X_07973__114 VPWR VGND net114 sg13g2_tiehi
X_06892_ VGND VPWR net1095 _02896_ _00691_ _02897_ sg13g2_a21oi_1
X_08631_ net1766 VGND VPWR net2636 i_exotiny._0029_\[0\] clknet_leaf_143_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_12_0 VPWR VGND sg13g2_fill_1
XFILLER_95_996 VPWR VGND sg13g2_decap_8
XFILLER_54_304 VPWR VGND sg13g2_fill_1
X_05843_ _02432_ _02431_ _02050_ _02051_ _01496_ VPWR VGND sg13g2_a22oi_1
X_05774_ _02400_ i_exotiny._2034_\[5\] _00026_ VPWR VGND sg13g2_nand2_1
X_08562_ net80 VGND VPWR net3518 i_exotiny._0314_\[7\] clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
XFILLER_35_540 VPWR VGND sg13g2_fill_1
X_08493_ net187 VGND VPWR net2877 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[13\]
+ clknet_leaf_71_clk_regs sg13g2_dfrbpq_1
X_07513_ net3377 net3113 net904 _01096_ VPWR VGND sg13g2_mux2_1
X_04725_ _01481_ VPWR _01482_ VGND _01380_ _01453_ sg13g2_o21ai_1
X_04656_ VPWR _01418_ net2 VGND sg13g2_inv_1
X_07444_ _03085_ VPWR _01055_ VGND net1081 _03084_ sg13g2_o21ai_1
X_08342__336 VPWR VGND net336 sg13g2_tiehi
X_07375_ net3584 net1213 _03032_ VPWR VGND sg13g2_and2_1
X_06326_ net2429 net1976 net1035 _00463_ VPWR VGND sg13g2_mux2_1
X_09114_ net868 VGND VPWR _01169_ i_exotiny._0030_\[2\] clknet_leaf_157_clk_regs sg13g2_dfrbpq_2
X_06257_ net2640 net3159 net1039 _00406_ VPWR VGND sg13g2_mux2_1
X_09045_ net1358 VGND VPWR _01102_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[0\]
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
Xclkbuf_leaf_19_clk_regs clknet_5_13__leaf_clk_regs clknet_leaf_19_clk_regs VPWR VGND
+ sg13g2_buf_8
X_05208_ _01936_ _01790_ i_exotiny._0034_\[1\] _01788_ i_exotiny._0039_\[1\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_104_523 VPWR VGND sg13g2_decap_8
XFILLER_89_212 VPWR VGND sg13g2_fill_1
X_06188_ _02539_ _01365_ net1105 VPWR VGND sg13g2_nand2_1
Xhold463 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[30\]
+ VPWR VGND net2290 sg13g2_dlygate4sd3_1
Xhold452 _00717_ VPWR VGND net2279 sg13g2_dlygate4sd3_1
XFILLER_2_628 VPWR VGND sg13g2_fill_1
Xhold430 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[24\]
+ VPWR VGND net2257 sg13g2_dlygate4sd3_1
Xhold441 _01324_ VPWR VGND net2268 sg13g2_dlygate4sd3_1
XFILLER_104_556 VPWR VGND sg13g2_decap_8
Xclkbuf_5_31__f_clk_regs clknet_4_15_0_clk_regs clknet_5_31__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold485 _00972_ VPWR VGND net2312 sg13g2_dlygate4sd3_1
Xhold496 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[16\]
+ VPWR VGND net2323 sg13g2_dlygate4sd3_1
Xhold474 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[9\]
+ VPWR VGND net2301 sg13g2_dlygate4sd3_1
X_05139_ VGND VPWR _01869_ _01868_ _01846_ sg13g2_or2_1
Xfanout910 net912 net910 VPWR VGND sg13g2_buf_8
Xfanout943 net944 net943 VPWR VGND sg13g2_buf_8
Xfanout932 _02621_ net932 VPWR VGND sg13g2_buf_8
Xfanout921 net922 net921 VPWR VGND sg13g2_buf_8
Xfanout976 net977 net976 VPWR VGND sg13g2_buf_8
Xfanout954 _02534_ net954 VPWR VGND sg13g2_buf_8
Xfanout965 _02511_ net965 VPWR VGND sg13g2_buf_8
XFILLER_85_440 VPWR VGND sg13g2_fill_1
Xhold1130 _00918_ VPWR VGND net2957 sg13g2_dlygate4sd3_1
Xhold1141 _00843_ VPWR VGND net2968 sg13g2_dlygate4sd3_1
Xfanout998 net999 net998 VPWR VGND sg13g2_buf_8
Xfanout987 _03223_ net987 VPWR VGND sg13g2_buf_8
X_08829_ net1579 VGND VPWR _00887_ i_exotiny.i_wb_spi.state_r\[28\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
Xhold1185 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[22\]
+ VPWR VGND net3012 sg13g2_dlygate4sd3_1
XFILLER_57_186 VPWR VGND sg13g2_fill_2
Xhold1163 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[8\]
+ VPWR VGND net2990 sg13g2_dlygate4sd3_1
Xhold1152 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[13\]
+ VPWR VGND net2979 sg13g2_dlygate4sd3_1
Xhold1174 _00831_ VPWR VGND net3001 sg13g2_dlygate4sd3_1
X_08034__660 VPWR VGND net660 sg13g2_tiehi
Xhold1196 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[29\]
+ VPWR VGND net3023 sg13g2_dlygate4sd3_1
XFILLER_72_145 VPWR VGND sg13g2_fill_1
XFILLER_57_197 VPWR VGND sg13g2_fill_2
XFILLER_14_735 VPWR VGND sg13g2_fill_2
XFILLER_13_245 VPWR VGND sg13g2_fill_2
XFILLER_10_963 VPWR VGND sg13g2_decap_8
Xclkload19 clkload19/Y clknet_leaf_9_clk_regs VPWR VGND sg13g2_inv_2
XFILLER_6_934 VPWR VGND sg13g2_decap_8
X_08041__653 VPWR VGND net653 sg13g2_tiehi
XFILLER_92_977 VPWR VGND sg13g2_decap_8
XFILLER_36_337 VPWR VGND sg13g2_fill_2
X_05490_ _02185_ VPWR i_exotiny._1611_\[10\] VGND net1074 _02187_ sg13g2_o21ai_1
X_07160_ net2213 net2198 net1008 _00908_ VPWR VGND sg13g2_mux2_1
X_07091_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[19\]
+ net2117 net914 _00846_ VPWR VGND sg13g2_mux2_1
X_06111_ _02518_ _02525_ _02526_ VPWR VGND sg13g2_nor2_2
X_06042_ net2563 net2766 net962 _00227_ VPWR VGND sg13g2_mux2_1
XFILLER_99_521 VPWR VGND sg13g2_decap_4
X_07993_ net134 VGND VPWR net3597 i_exotiny._0369_\[3\] clknet_leaf_15_clk_regs sg13g2_dfrbpq_2
XFILLER_55_602 VPWR VGND sg13g2_decap_4
X_06944_ net2192 net2734 net926 _00723_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_137_clk_regs clknet_5_21__leaf_clk_regs clknet_leaf_137_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_95_782 VPWR VGND sg13g2_fill_2
XFILLER_94_270 VPWR VGND sg13g2_decap_8
X_06875_ net3601 net1189 _02883_ VPWR VGND sg13g2_nor2_1
X_05826_ net2504 net2247 net1054 _00098_ VPWR VGND sg13g2_mux2_1
X_08614_ net1782 VGND VPWR net3615 i_exotiny._1616_\[2\] clknet_leaf_23_clk_regs sg13g2_dfrbpq_2
X_08485__195 VPWR VGND net195 sg13g2_tiehi
X_08545_ net111 VGND VPWR net3758 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[1\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_2
X_05757_ _02389_ _02388_ net1991 _02367_ _01577_ VPWR VGND sg13g2_a22oi_1
X_05688_ net1122 net1926 _02337_ VPWR VGND sg13g2_nor2b_1
X_08476_ net204 VGND VPWR net3329 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[28\]
+ clknet_leaf_115_clk_regs sg13g2_dfrbpq_1
XFILLER_24_36 VPWR VGND sg13g2_fill_2
X_04708_ net1253 _01457_ _01466_ VPWR VGND sg13g2_and2_1
X_04639_ VPWR _01401_ i_exotiny._2034_\[3\] VGND sg13g2_inv_1
X_07427_ net1081 net2040 _03072_ _01051_ VPWR VGND sg13g2_a21o_1
X_07358_ _03019_ _03009_ _03018_ net1207 net1949 VPWR VGND sg13g2_a22oi_1
X_06309_ net3263 net3044 net1033 _00446_ VPWR VGND sg13g2_mux2_1
X_07289_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[14\]
+ net2035 net909 _01006_ VPWR VGND sg13g2_mux2_1
X_09028_ net1374 VGND VPWR net3662 i_exotiny._0315_\[16\] clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
XFILLER_105_832 VPWR VGND sg13g2_decap_8
XFILLER_104_320 VPWR VGND sg13g2_decap_8
Xhold260 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.genblk7.g_value.r_value[0]
+ VPWR VGND net2087 sg13g2_dlygate4sd3_1
X_08492__188 VPWR VGND net188 sg13g2_tiehi
Xhold271 _01139_ VPWR VGND net2098 sg13g2_dlygate4sd3_1
X_08318__360 VPWR VGND net360 sg13g2_tiehi
Xhold282 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[20\]
+ VPWR VGND net2109 sg13g2_dlygate4sd3_1
Xhold293 _00412_ VPWR VGND net2120 sg13g2_dlygate4sd3_1
XFILLER_104_397 VPWR VGND sg13g2_decap_8
XFILLER_46_613 VPWR VGND sg13g2_fill_2
XFILLER_74_999 VPWR VGND sg13g2_fill_2
XFILLER_92_1012 VPWR VGND sg13g2_decap_8
X_08325__353 VPWR VGND net353 sg13g2_tiehi
XFILLER_5_241 VPWR VGND sg13g2_fill_2
XFILLER_96_502 VPWR VGND sg13g2_fill_1
XFILLER_69_727 VPWR VGND sg13g2_fill_1
XFILLER_2_992 VPWR VGND sg13g2_decap_8
X_08332__346 VPWR VGND net346 sg13g2_tiehi
X_04990_ _01721_ _01707_ _01722_ VPWR VGND _01717_ sg13g2_nand3b_1
Xinput6 ui_in[4] net6 VPWR VGND sg13g2_buf_1
XFILLER_77_782 VPWR VGND sg13g2_fill_1
XFILLER_37_602 VPWR VGND sg13g2_fill_1
X_06660_ net1162 VPWR _02700_ VGND i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data[0]
+ _02691_ sg13g2_o21ai_1
X_05611_ net1907 net1061 _02279_ VPWR VGND sg13g2_nor2_1
X_06591_ net1199 _02649_ _02650_ _00637_ VPWR VGND sg13g2_nor3_1
X_08330_ net348 VGND VPWR net3180 i_exotiny._0016_\[0\] clknet_leaf_99_clk_regs sg13g2_dfrbpq_2
X_05542_ net1277 net3549 _02228_ VPWR VGND sg13g2_nor2b_1
X_09191__790 VPWR VGND net790 sg13g2_tiehi
X_08261_ net416 VGND VPWR _00342_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[28\]
+ clknet_leaf_56_clk_regs sg13g2_dfrbpq_1
X_05473_ net1265 i_exotiny._1711_ _01521_ _02175_ VPWR VGND sg13g2_nor3_1
X_07212_ VGND VPWR _01415_ net1088 _00941_ _02967_ sg13g2_a21oi_1
X_08192_ net485 VGND VPWR net2436 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[23\]
+ clknet_leaf_69_clk_regs sg13g2_dfrbpq_1
X_07143_ net2174 i_exotiny._0036_\[0\] net1011 _00891_ VPWR VGND sg13g2_mux2_1
XFILLER_106_629 VPWR VGND sg13g2_decap_8
X_08024__670 VPWR VGND net670 sg13g2_tiehi
X_07074_ net3080 net3073 net916 _00829_ VPWR VGND sg13g2_mux2_1
X_06025_ _00022_ net1103 _02507_ VPWR VGND sg13g2_nor2_1
X_07979__120 VPWR VGND net120 sg13g2_tiehi
XFILLER_102_846 VPWR VGND sg13g2_decap_8
XFILLER_99_395 VPWR VGND sg13g2_decap_8
XFILLER_101_345 VPWR VGND sg13g2_decap_8
X_07976_ net117 VGND VPWR net3595 i_exotiny._0369_\[29\] clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
X_08844__1142 VPWR VGND net1562 sg13g2_tiehi
X_06927_ net2721 net2848 net927 _00706_ VPWR VGND sg13g2_mux2_1
XFILLER_67_281 VPWR VGND sg13g2_fill_2
XFILLER_16_808 VPWR VGND sg13g2_decap_4
X_06858_ net1171 VPWR _02869_ VGND i_exotiny.i_wb_spi.dat_rx_r\[26\] net1186 sg13g2_o21ai_1
X_08031__663 VPWR VGND net663 sg13g2_tiehi
X_05809_ net2815 i_exotiny._0018_\[1\] net1056 _00081_ VPWR VGND sg13g2_mux2_1
X_06789_ net3596 net1188 _02811_ VPWR VGND sg13g2_nor2_1
XFILLER_27_178 VPWR VGND sg13g2_fill_2
X_08528_ net152 VGND VPWR net2702 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[16\]
+ clknet_leaf_176_clk_regs sg13g2_dfrbpq_1
X_08459_ net221 VGND VPWR _00533_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[11\]
+ clknet_leaf_159_clk_regs sg13g2_dfrbpq_1
Xclkbuf_leaf_34_clk_regs clknet_5_9__leaf_clk_regs clknet_leaf_34_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_51_34 VPWR VGND sg13g2_fill_1
XFILLER_3_767 VPWR VGND sg13g2_decap_8
XFILLER_104_194 VPWR VGND sg13g2_decap_8
XFILLER_78_568 VPWR VGND sg13g2_fill_2
XFILLER_76_42 VPWR VGND sg13g2_fill_1
X_08795__1193 VPWR VGND net1613 sg13g2_tiehi
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_74_774 VPWR VGND sg13g2_fill_2
XFILLER_62_914 VPWR VGND sg13g2_fill_2
XFILLER_18_145 VPWR VGND sg13g2_fill_2
XFILLER_46_498 VPWR VGND sg13g2_fill_1
XFILLER_41_181 VPWR VGND sg13g2_fill_1
XFILLER_42_693 VPWR VGND sg13g2_decap_8
XFILLER_30_888 VPWR VGND sg13g2_fill_1
X_08008__687 VPWR VGND net687 sg13g2_tiehi
XFILLER_97_877 VPWR VGND sg13g2_decap_8
XFILLER_96_343 VPWR VGND sg13g2_decap_8
XFILLER_57_719 VPWR VGND sg13g2_fill_1
Xhold1707 _00919_ VPWR VGND net3534 sg13g2_dlygate4sd3_1
X_07830_ net3048 net2162 net984 _01303_ VPWR VGND sg13g2_mux2_1
X_07761_ net2241 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[13\]
+ net992 _01246_ VPWR VGND sg13g2_mux2_1
Xhold1729 i_exotiny.i_wb_spi.dat_rx_r\[3\] VPWR VGND net3556 sg13g2_dlygate4sd3_1
XFILLER_2_50 VPWR VGND sg13g2_fill_1
Xhold1718 i_exotiny._0315_\[13\] VPWR VGND net3545 sg13g2_dlygate4sd3_1
X_09078__904 VPWR VGND net1324 sg13g2_tiehi
X_06712_ i_exotiny._0369_\[3\] i_exotiny.i_wb_spi.dat_rx_r\[3\] net1193 _02746_ VPWR
+ VGND sg13g2_mux2_1
X_04973_ _01705_ _01393_ _01703_ VPWR VGND sg13g2_xnor2_1
X_07692_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[27\]
+ net2209 net999 _01194_ VPWR VGND sg13g2_mux2_1
XFILLER_37_454 VPWR VGND sg13g2_fill_2
XFILLER_64_262 VPWR VGND sg13g2_fill_1
X_06643_ net1974 net1161 _02685_ VPWR VGND sg13g2_nor2_1
X_09256__551 VPWR VGND net551 sg13g2_tiehi
X_06574_ i_exotiny._0314_\[4\] net1160 _02639_ VPWR VGND sg13g2_nor2_1
X_08313_ net365 VGND VPWR _00394_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[15\]
+ clknet_leaf_74_clk_regs sg13g2_dfrbpq_1
X_08482__198 VPWR VGND net198 sg13g2_tiehi
X_05525_ VGND VPWR i_exotiny._0314_\[14\] net1276 _02214_ _02213_ sg13g2_a21oi_1
X_08308__370 VPWR VGND net370 sg13g2_tiehi
X_09293_ net1813 VGND VPWR _01348_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[19\]
+ clknet_leaf_167_clk_regs sg13g2_dfrbpq_1
X_08244_ net433 VGND VPWR net2740 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[11\]
+ clknet_leaf_60_clk_regs sg13g2_dfrbpq_1
X_05456_ _02163_ _02146_ i_exotiny._1616_\[2\] _02145_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data[0]
+ VPWR VGND sg13g2_a22oi_1
X_05387_ VGND VPWR _02094_ _02106_ _02107_ _02096_ sg13g2_a21oi_1
X_08175_ net502 VGND VPWR _00256_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[6\]
+ clknet_leaf_70_clk_regs sg13g2_dfrbpq_1
X_07126_ net1290 net1859 _00876_ VPWR VGND sg13g2_and2_1
XFILLER_106_426 VPWR VGND sg13g2_decap_8
X_07057_ net2555 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[23\]
+ net1016 _00818_ VPWR VGND sg13g2_mux2_1
XFILLER_82_1011 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_152_clk_regs clknet_5_18__leaf_clk_regs clknet_leaf_152_clk_regs VPWR
+ VGND sg13g2_buf_8
X_06008_ net2758 net873 _02493_ _02498_ VPWR VGND sg13g2_mux2_1
X_08315__363 VPWR VGND net363 sg13g2_tiehi
XFILLER_29_922 VPWR VGND sg13g2_fill_2
X_07959_ net1176 VGND VPWR net3736 i_exotiny.i_wdg_top.o_wb_dat\[0\] clknet_leaf_37_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_56_752 VPWR VGND sg13g2_fill_1
XFILLER_29_977 VPWR VGND sg13g2_fill_2
XFILLER_70_210 VPWR VGND sg13g2_fill_1
XFILLER_43_457 VPWR VGND sg13g2_fill_2
XFILLER_70_298 VPWR VGND sg13g2_fill_2
XFILLER_11_332 VPWR VGND sg13g2_fill_1
XFILLER_8_804 VPWR VGND sg13g2_fill_1
X_08322__356 VPWR VGND net356 sg13g2_tiehi
X_08703__1285 VPWR VGND net1705 sg13g2_tiehi
XFILLER_106_993 VPWR VGND sg13g2_decap_8
XFILLER_3_586 VPWR VGND sg13g2_fill_1
XFILLER_66_505 VPWR VGND sg13g2_fill_1
X_08925__1057 VPWR VGND net1477 sg13g2_tiehi
XFILLER_47_752 VPWR VGND sg13g2_fill_1
XFILLER_46_240 VPWR VGND sg13g2_fill_1
X_08014__680 VPWR VGND net680 sg13g2_tiehi
XFILLER_61_243 VPWR VGND sg13g2_fill_1
X_06290_ net3229 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[22\]
+ net941 _00433_ VPWR VGND sg13g2_mux2_1
X_05310_ i_exotiny._0036_\[0\] _01644_ _02036_ VPWR VGND sg13g2_nor2_1
X_05241_ VGND VPWR i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[1\].i_hadd.a_i
+ _01612_ _01969_ _01968_ sg13g2_a21oi_1
X_05172_ net1110 _01897_ _01901_ VPWR VGND sg13g2_nor2_1
XFILLER_6_380 VPWR VGND sg13g2_fill_2
Xhold826 _00899_ VPWR VGND net2653 sg13g2_dlygate4sd3_1
Xhold815 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[22\]
+ VPWR VGND net2642 sg13g2_dlygate4sd3_1
Xhold837 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[30\]
+ VPWR VGND net2664 sg13g2_dlygate4sd3_1
Xhold804 _00203_ VPWR VGND net2631 sg13g2_dlygate4sd3_1
Xhold848 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[4\]
+ VPWR VGND net2675 sg13g2_dlygate4sd3_1
Xhold859 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[10\]
+ VPWR VGND net2686 sg13g2_dlygate4sd3_1
XFILLER_42_0 VPWR VGND sg13g2_fill_2
X_08021__673 VPWR VGND net673 sg13g2_tiehi
X_08931_ net1471 VGND VPWR net2399 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[29\]
+ clknet_leaf_113_clk_regs sg13g2_dfrbpq_1
X_08862_ net1544 VGND VPWR net2661 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[29\]
+ clknet_leaf_186_clk_regs sg13g2_dfrbpq_1
Xhold1526 _00975_ VPWR VGND net3353 sg13g2_dlygate4sd3_1
Xhold1515 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[26\]
+ VPWR VGND net3342 sg13g2_dlygate4sd3_1
X_07813_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[27\]
+ net2497 net891 _01292_ VPWR VGND sg13g2_mux2_1
Xhold1504 _00842_ VPWR VGND net3331 sg13g2_dlygate4sd3_1
Xhold1559 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[11\]
+ VPWR VGND net3386 sg13g2_dlygate4sd3_1
Xhold1548 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[29\]
+ VPWR VGND net3375 sg13g2_dlygate4sd3_1
X_08793_ net1615 VGND VPWR net2695 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[24\]
+ clknet_leaf_167_clk_regs sg13g2_dfrbpq_1
Xhold1537 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[14\]
+ VPWR VGND net3364 sg13g2_dlygate4sd3_1
X_07744_ net1116 net1060 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data[0]
+ _03209_ VPWR VGND sg13g2_nand3_1
X_04956_ _01688_ _01425_ _01687_ VPWR VGND sg13g2_xnor2_1
XFILLER_93_880 VPWR VGND sg13g2_fill_1
X_07675_ net3062 net3434 net1002 _01177_ VPWR VGND sg13g2_mux2_1
X_04887_ i_exotiny._0077_\[2\] i_exotiny._0077_\[3\] net1255 _01619_ VGND VPWR _01613_
+ sg13g2_nor4_2
XFILLER_13_608 VPWR VGND sg13g2_fill_1
X_06626_ net2008 net1152 _02674_ VPWR VGND sg13g2_nor2_1
XFILLER_40_438 VPWR VGND sg13g2_fill_1
X_06557_ net3787 net1259 net1211 _00624_ VPWR VGND sg13g2_mux2_1
X_06488_ net2940 net3195 net1023 _00569_ VPWR VGND sg13g2_mux2_1
X_09276_ net69 VGND VPWR net2452 i_exotiny._0021_\[2\] clknet_leaf_170_clk_regs sg13g2_dfrbpq_2
X_05508_ net1275 i_exotiny._0315_\[9\] _02201_ VPWR VGND sg13g2_nor2b_1
X_05439_ net1232 _02133_ _02142_ _02148_ VPWR VGND sg13g2_nor3_1
X_08227_ net450 VGND VPWR _00308_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[26\]
+ clknet_leaf_169_clk_regs sg13g2_dfrbpq_1
XFILLER_10_1005 VPWR VGND sg13g2_decap_8
XFILLER_106_223 VPWR VGND sg13g2_decap_8
X_08158_ net520 VGND VPWR net2700 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[22\]
+ clknet_leaf_133_clk_regs sg13g2_dfrbpq_1
X_08089_ net605 VGND VPWR _00170_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[26\]
+ clknet_leaf_85_clk_regs sg13g2_dfrbpq_1
X_07109_ VGND VPWR _01379_ _01579_ _00859_ _02946_ sg13g2_a21oi_1
XFILLER_103_930 VPWR VGND sg13g2_decap_8
XFILLER_0_556 VPWR VGND sg13g2_fill_1
XFILLER_102_462 VPWR VGND sg13g2_decap_8
XFILLER_87_173 VPWR VGND sg13g2_fill_2
XFILLER_44_700 VPWR VGND sg13g2_decap_8
XFILLER_56_593 VPWR VGND sg13g2_fill_1
XFILLER_16_413 VPWR VGND sg13g2_fill_2
X_08581__1400 VPWR VGND net1820 sg13g2_tiehi
XFILLER_16_479 VPWR VGND sg13g2_fill_2
XFILLER_106_1000 VPWR VGND sg13g2_decap_8
X_09068__914 VPWR VGND net1334 sg13g2_tiehi
XFILLER_4_862 VPWR VGND sg13g2_decap_8
X_09246__561 VPWR VGND net561 sg13g2_tiehi
XFILLER_106_790 VPWR VGND sg13g2_decap_8
Xfanout1140 net1141 net1140 VPWR VGND sg13g2_buf_1
Xfanout1173 _01516_ net1173 VPWR VGND sg13g2_buf_8
Xfanout1162 net1164 net1162 VPWR VGND sg13g2_buf_8
Xfanout1151 _02984_ net1151 VPWR VGND sg13g2_buf_2
X_05790_ _02410_ VPWR _00076_ VGND net1888 _01551_ sg13g2_o21ai_1
Xfanout1195 net1197 net1195 VPWR VGND sg13g2_buf_8
Xfanout1184 _01472_ net1184 VPWR VGND sg13g2_buf_8
X_04810_ VPWR VGND _01522_ _01553_ _01520_ net1265 _01554_ _01511_ sg13g2_a221oi_1
XFILLER_93_187 VPWR VGND sg13g2_fill_2
X_04741_ net1197 net1894 _00002_ VPWR VGND sg13g2_nor2_1
X_09075__907 VPWR VGND net1327 sg13g2_tiehi
XFILLER_23_939 VPWR VGND sg13g2_fill_1
XFILLER_35_788 VPWR VGND sg13g2_fill_2
X_04672_ net1248 net1250 net1252 _01433_ VGND VPWR net1253 sg13g2_nor4_2
X_07460_ _03096_ VPWR _01060_ VGND net1080 _03095_ sg13g2_o21ai_1
X_06411_ _01390_ net1233 i_exotiny._0315_\[4\] _02593_ VPWR VGND sg13g2_nor3_2
X_09253__554 VPWR VGND net554 sg13g2_tiehi
X_07391_ net3828 net1215 _03044_ VPWR VGND sg13g2_and2_1
X_06342_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[1\] _02474_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[2\]
+ _02564_ VPWR VGND sg13g2_nand3_1
X_09130_ net852 VGND VPWR _01185_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[18\]
+ clknet_leaf_156_clk_regs sg13g2_dfrbpq_1
X_09061_ net1341 VGND VPWR _01116_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[1\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_31_994 VPWR VGND sg13g2_fill_2
X_08305__373 VPWR VGND net373 sg13g2_tiehi
X_06273_ net2881 net2119 net939 _00416_ VPWR VGND sg13g2_mux2_1
X_08012_ net682 VGND VPWR _00093_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[13\]
+ clknet_leaf_69_clk_regs sg13g2_dfrbpq_1
Xhold612 _00992_ VPWR VGND net2439 sg13g2_dlygate4sd3_1
Xhold601 _00357_ VPWR VGND net2428 sg13g2_dlygate4sd3_1
X_05224_ _01952_ _01651_ i_exotiny._0039_\[1\] _01621_ i_exotiny._0043_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold634 _01240_ VPWR VGND net2461 sg13g2_dlygate4sd3_1
Xhold623 i_exotiny._0034_\[0\] VPWR VGND net2450 sg13g2_dlygate4sd3_1
Xhold645 _01325_ VPWR VGND net2472 sg13g2_dlygate4sd3_1
X_05155_ _01885_ _01649_ i_exotiny._0042_\[2\] _01647_ i_exotiny._0032_\[2\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_104_727 VPWR VGND sg13g2_decap_8
Xhold678 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[31\]
+ VPWR VGND net2505 sg13g2_dlygate4sd3_1
Xclkbuf_5_30__f_clk_regs clknet_4_15_0_clk_regs clknet_5_30__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold667 _00491_ VPWR VGND net2494 sg13g2_dlygate4sd3_1
Xhold656 _00112_ VPWR VGND net2483 sg13g2_dlygate4sd3_1
X_05086_ net1243 _01603_ _01817_ VPWR VGND sg13g2_nor2_1
XFILLER_103_248 VPWR VGND sg13g2_decap_8
Xhold689 _00498_ VPWR VGND net2516 sg13g2_dlygate4sd3_1
X_08914_ net1488 VGND VPWR net2312 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[12\]
+ clknet_leaf_65_clk_regs sg13g2_dfrbpq_1
Xhold2002 _02582_ VPWR VGND net3829 sg13g2_dlygate4sd3_1
XFILLER_98_972 VPWR VGND sg13g2_decap_8
XFILLER_97_471 VPWR VGND sg13g2_fill_2
XFILLER_57_302 VPWR VGND sg13g2_fill_1
Xhold2013 i_exotiny._1308_ VPWR VGND net3840 sg13g2_dlygate4sd3_1
XFILLER_97_482 VPWR VGND sg13g2_decap_8
Xhold1334 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[30\]
+ VPWR VGND net3161 sg13g2_dlygate4sd3_1
Xhold1301 _00314_ VPWR VGND net3128 sg13g2_dlygate4sd3_1
Xhold1323 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[26\]
+ VPWR VGND net3150 sg13g2_dlygate4sd3_1
X_08845_ net1561 VGND VPWR net2324 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[12\]
+ clknet_leaf_185_clk_regs sg13g2_dfrbpq_1
Xhold1312 _01180_ VPWR VGND net3139 sg13g2_dlygate4sd3_1
XFILLER_100_966 VPWR VGND sg13g2_decap_8
X_08312__366 VPWR VGND net366 sg13g2_tiehi
Xhold1367 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[14\]
+ VPWR VGND net3194 sg13g2_dlygate4sd3_1
XFILLER_85_677 VPWR VGND sg13g2_fill_2
XFILLER_57_346 VPWR VGND sg13g2_fill_1
X_08776_ net1632 VGND VPWR _00834_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[7\]
+ clknet_leaf_164_clk_regs sg13g2_dfrbpq_1
Xhold1345 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[25\]
+ VPWR VGND net3172 sg13g2_dlygate4sd3_1
Xhold1356 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[27\]
+ VPWR VGND net3183 sg13g2_dlygate4sd3_1
Xhold1378 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[12\]
+ VPWR VGND net3205 sg13g2_dlygate4sd3_1
Xhold1389 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[14\]
+ VPWR VGND net3216 sg13g2_dlygate4sd3_1
XFILLER_57_379 VPWR VGND sg13g2_fill_2
X_05988_ net2377 net3296 net1048 _00190_ VPWR VGND sg13g2_mux2_1
X_07727_ net2839 net2048 net993 _01223_ VPWR VGND sg13g2_mux2_1
X_04939_ VPWR VGND i_exotiny._0039_\[3\] _01670_ _01651_ i_exotiny._0032_\[3\] _01671_
+ _01647_ sg13g2_a221oi_1
X_07658_ net2888 _03190_ net898 _01164_ VPWR VGND sg13g2_mux2_1
X_07589_ net2028 _03163_ _03164_ VPWR VGND sg13g2_nor2_1
X_06609_ net1198 _02661_ _02662_ _00643_ VPWR VGND sg13g2_nor3_1
X_09259_ net243 VGND VPWR _01314_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[17\]
+ clknet_leaf_128_clk_regs sg13g2_dfrbpq_1
XFILLER_1_810 VPWR VGND sg13g2_decap_8
XFILLER_68_32 VPWR VGND sg13g2_fill_1
XFILLER_76_611 VPWR VGND sg13g2_fill_2
XFILLER_1_887 VPWR VGND sg13g2_decap_8
XFILLER_64_817 VPWR VGND sg13g2_fill_1
XFILLER_95_1010 VPWR VGND sg13g2_decap_8
Xhold1890 i_exotiny._1617_\[0\] VPWR VGND net3717 sg13g2_dlygate4sd3_1
XFILLER_31_224 VPWR VGND sg13g2_fill_1
XFILLER_9_932 VPWR VGND sg13g2_decap_8
XFILLER_13_983 VPWR VGND sg13g2_decap_8
XFILLER_99_736 VPWR VGND sg13g2_fill_1
XFILLER_98_202 VPWR VGND sg13g2_fill_1
XFILLER_99_747 VPWR VGND sg13g2_fill_2
XFILLER_98_257 VPWR VGND sg13g2_decap_8
XFILLER_67_600 VPWR VGND sg13g2_fill_2
X_06960_ i_exotiny._0034_\[2\] net2243 net1022 _00733_ VPWR VGND sg13g2_mux2_1
X_05911_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[16\]
+ net2357 net976 _00128_ VPWR VGND sg13g2_mux2_1
X_06891_ net3747 net1095 _02897_ VPWR VGND sg13g2_nor2_1
XFILLER_95_975 VPWR VGND sg13g2_decap_8
X_08630_ net1768 VGND VPWR i_exotiny._1489_\[3\] i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[3\]
+ clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
X_05842_ _01496_ _01497_ _02431_ VPWR VGND sg13g2_nor2_2
X_05773_ _02399_ VPWR _00070_ VGND net1143 _02398_ sg13g2_o21ai_1
X_08561_ net82 VGND VPWR _00634_ i_exotiny._0314_\[6\] clknet_leaf_166_clk_regs sg13g2_dfrbpq_1
X_08492_ net188 VGND VPWR _00566_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[12\]
+ clknet_leaf_108_clk_regs sg13g2_dfrbpq_1
X_07512_ i_exotiny._0315_\[29\] net3220 net901 _01095_ VPWR VGND sg13g2_mux2_1
X_04724_ i_exotiny._1265_ _01464_ net1268 _01481_ VPWR VGND sg13g2_nand3_1
XFILLER_90_680 VPWR VGND sg13g2_fill_2
X_04655_ _01417_ i_exotiny.i_wb_spi.dat_rx_r\[17\] VPWR VGND sg13g2_inv_2
X_07443_ VGND VPWR net3565 net1081 _03085_ _03077_ sg13g2_a21oi_1
X_09113_ net869 VGND VPWR _01168_ i_exotiny._0030_\[1\] clknet_leaf_154_clk_regs sg13g2_dfrbpq_2
X_07374_ net1949 net1077 _03031_ VPWR VGND sg13g2_nor2_1
X_06325_ net2000 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[19\]
+ net1036 _00462_ VPWR VGND sg13g2_mux2_1
X_06256_ net3136 net2915 net1038 _00405_ VPWR VGND sg13g2_mux2_1
X_09044_ net1359 VGND VPWR i_exotiny._1206_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r
+ clknet_5_2__leaf_clk_regs sg13g2_dfrbpq_1
Xhold420 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[18\]
+ VPWR VGND net2247 sg13g2_dlygate4sd3_1
X_05207_ _01935_ _01791_ i_exotiny._0026_\[1\] _01785_ i_exotiny._0043_\[1\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_104_502 VPWR VGND sg13g2_decap_8
Xhold442 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[11\]
+ VPWR VGND net2269 sg13g2_dlygate4sd3_1
X_06187_ net3174 _02538_ net950 _00345_ VPWR VGND sg13g2_mux2_1
X_08920__1062 VPWR VGND net1482 sg13g2_tiehi
Xhold453 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[19\]
+ VPWR VGND net2280 sg13g2_dlygate4sd3_1
Xhold431 _00237_ VPWR VGND net2258 sg13g2_dlygate4sd3_1
XFILLER_104_546 VPWR VGND sg13g2_fill_1
Xhold486 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[30\]
+ VPWR VGND net2313 sg13g2_dlygate4sd3_1
Xhold464 _01018_ VPWR VGND net2291 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_59_clk_regs clknet_5_12__leaf_clk_regs clknet_leaf_59_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold475 _01176_ VPWR VGND net2302 sg13g2_dlygate4sd3_1
Xfanout900 _03188_ net900 VPWR VGND sg13g2_buf_8
X_05138_ _01855_ _01858_ _01867_ _01868_ VPWR VGND sg13g2_nor3_2
Xfanout911 net912 net911 VPWR VGND sg13g2_buf_8
Xfanout933 _02621_ net933 VPWR VGND sg13g2_buf_1
Xhold497 _00903_ VPWR VGND net2324 sg13g2_dlygate4sd3_1
Xfanout922 net923 net922 VPWR VGND sg13g2_buf_8
X_05069_ _01794_ _01795_ _01775_ _01801_ VPWR VGND _01800_ sg13g2_nand4_1
Xfanout966 net971 net966 VPWR VGND sg13g2_buf_8
Xfanout977 _02479_ net977 VPWR VGND sg13g2_buf_8
Xfanout944 _02553_ net944 VPWR VGND sg13g2_buf_8
Xfanout955 net956 net955 VPWR VGND sg13g2_buf_8
Xhold1142 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[14\]
+ VPWR VGND net2969 sg13g2_dlygate4sd3_1
Xfanout988 _03211_ net988 VPWR VGND sg13g2_buf_8
XFILLER_86_964 VPWR VGND sg13g2_fill_2
Xhold1120 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[9\]
+ VPWR VGND net2947 sg13g2_dlygate4sd3_1
Xhold1131 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[12\]
+ VPWR VGND net2958 sg13g2_dlygate4sd3_1
Xfanout999 _03194_ net999 VPWR VGND sg13g2_buf_8
X_08828_ net1580 VGND VPWR _00886_ i_exotiny.i_wb_spi.state_r\[27\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_86_997 VPWR VGND sg13g2_decap_8
XFILLER_58_688 VPWR VGND sg13g2_fill_1
XFILLER_57_176 VPWR VGND sg13g2_fill_1
XFILLER_57_154 VPWR VGND sg13g2_fill_1
Xhold1164 _01203_ VPWR VGND net2991 sg13g2_dlygate4sd3_1
Xhold1153 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[8\]
+ VPWR VGND net2980 sg13g2_dlygate4sd3_1
Xhold1175 i_exotiny._0015_\[3\] VPWR VGND net3002 sg13g2_dlygate4sd3_1
X_08626__741 VPWR VGND net741 sg13g2_tiehi
Xhold1186 i_exotiny._0042_\[3\] VPWR VGND net3013 sg13g2_dlygate4sd3_1
X_08759_ net1649 VGND VPWR net3276 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[22\]
+ clknet_leaf_84_clk_regs sg13g2_dfrbpq_1
Xhold1197 _00343_ VPWR VGND net3024 sg13g2_dlygate4sd3_1
XFILLER_38_390 VPWR VGND sg13g2_fill_2
XFILLER_60_319 VPWR VGND sg13g2_fill_1
X_09058__924 VPWR VGND net1344 sg13g2_tiehi
XFILLER_54_861 VPWR VGND sg13g2_fill_2
XFILLER_53_393 VPWR VGND sg13g2_fill_2
XFILLER_26_585 VPWR VGND sg13g2_fill_1
XFILLER_16_1011 VPWR VGND sg13g2_fill_2
XFILLER_103_1014 VPWR VGND sg13g2_decap_8
XFILLER_10_942 VPWR VGND sg13g2_decap_8
XFILLER_70_88 VPWR VGND sg13g2_fill_1
XFILLER_6_913 VPWR VGND sg13g2_decap_8
X_09065__917 VPWR VGND net1337 sg13g2_tiehi
X_07996__137 VPWR VGND net137 sg13g2_tiehi
X_08740__1248 VPWR VGND net1668 sg13g2_tiehi
X_09243__564 VPWR VGND net564 sg13g2_tiehi
XFILLER_76_452 VPWR VGND sg13g2_fill_2
XFILLER_92_956 VPWR VGND sg13g2_decap_8
XFILLER_63_168 VPWR VGND sg13g2_fill_2
XFILLER_17_552 VPWR VGND sg13g2_fill_1
X_09250__557 VPWR VGND net557 sg13g2_tiehi
X_06110_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[1\] _02418_ _02525_
+ VPWR VGND net1262 sg13g2_nand3b_1
X_07090_ net3367 net3440 net917 _00845_ VPWR VGND sg13g2_mux2_1
X_08302__376 VPWR VGND net376 sg13g2_tiehi
X_06041_ net2604 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[9\]
+ net961 _00226_ VPWR VGND sg13g2_mux2_1
XFILLER_99_500 VPWR VGND sg13g2_decap_8
XFILLER_87_717 VPWR VGND sg13g2_fill_1
X_07992_ net133 VGND VPWR i_exotiny._1611_\[26\] i_exotiny._0369_\[2\] clknet_leaf_166_clk_regs
+ sg13g2_dfrbpq_2
X_08716__1272 VPWR VGND net1692 sg13g2_tiehi
X_06943_ net2315 net2488 net927 _00722_ VPWR VGND sg13g2_mux2_1
XFILLER_68_975 VPWR VGND sg13g2_fill_1
XFILLER_95_772 VPWR VGND sg13g2_fill_1
X_06874_ VGND VPWR net1094 _02881_ _00688_ _02882_ sg13g2_a21oi_1
X_05825_ net2543 net2745 net1057 _00097_ VPWR VGND sg13g2_mux2_1
X_08611__1365 VPWR VGND net1785 sg13g2_tiehi
X_08613_ net1783 VGND VPWR net3573 i_exotiny._1616_\[1\] clknet_leaf_22_clk_regs sg13g2_dfrbpq_2
X_05756_ VGND VPWR net3400 _02388_ _00064_ _01580_ sg13g2_a21oi_1
XFILLER_54_146 VPWR VGND sg13g2_fill_2
X_08544_ net112 VGND VPWR net3592 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[0\]
+ clknet_leaf_18_clk_regs sg13g2_dfrbpq_1
Xclkbuf_leaf_177_clk_regs clknet_5_1__leaf_clk_regs clknet_leaf_177_clk_regs VPWR
+ VGND sg13g2_buf_8
Xclkbuf_leaf_106_clk_regs clknet_5_28__leaf_clk_regs clknet_leaf_106_clk_regs VPWR
+ VGND sg13g2_buf_8
X_04707_ _01462_ _01463_ net1249 _01465_ VPWR VGND sg13g2_nand3_1
X_08938__1044 VPWR VGND net1464 sg13g2_tiehi
X_05687_ net2046 net1064 _02336_ VPWR VGND sg13g2_nor2_1
XFILLER_24_48 VPWR VGND sg13g2_fill_1
X_08475_ net205 VGND VPWR _00549_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[27\]
+ clknet_leaf_158_clk_regs sg13g2_dfrbpq_1
X_04638_ VPWR _01400_ i_exotiny._2034_\[2\] VGND sg13g2_inv_1
XFILLER_11_728 VPWR VGND sg13g2_fill_2
X_07426_ net1081 _03070_ _03071_ _03072_ VPWR VGND sg13g2_nor3_1
X_07357_ net2061 net1214 _03018_ VPWR VGND sg13g2_and2_1
X_06308_ net3519 net3674 net1037 _00445_ VPWR VGND sg13g2_mux2_1
X_07288_ net2067 net2127 net908 _01005_ VPWR VGND sg13g2_mux2_1
X_09027_ net1375 VGND VPWR net3613 i_exotiny._0315_\[15\] clknet_leaf_179_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_105_811 VPWR VGND sg13g2_decap_8
X_06239_ net3211 net2416 net1040 _00388_ VPWR VGND sg13g2_mux2_1
XFILLER_85_1020 VPWR VGND sg13g2_decap_8
Xhold261 _00346_ VPWR VGND net2088 sg13g2_dlygate4sd3_1
XFILLER_3_949 VPWR VGND sg13g2_decap_8
Xhold250 i_exotiny._1160_\[12\] VPWR VGND net2077 sg13g2_dlygate4sd3_1
XFILLER_105_888 VPWR VGND sg13g2_decap_8
Xhold283 _00330_ VPWR VGND net2110 sg13g2_dlygate4sd3_1
Xhold272 i_exotiny._0315_\[28\] VPWR VGND net2099 sg13g2_dlygate4sd3_1
Xhold294 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[30\]
+ VPWR VGND net2121 sg13g2_dlygate4sd3_1
XFILLER_104_376 VPWR VGND sg13g2_decap_8
XFILLER_77_238 VPWR VGND sg13g2_fill_1
XFILLER_85_260 VPWR VGND sg13g2_fill_1
XFILLER_19_817 VPWR VGND sg13g2_fill_2
XFILLER_45_102 VPWR VGND sg13g2_fill_2
XFILLER_74_967 VPWR VGND sg13g2_fill_1
XFILLER_14_511 VPWR VGND sg13g2_fill_1
XFILLER_26_360 VPWR VGND sg13g2_fill_2
XFILLER_60_138 VPWR VGND sg13g2_fill_1
X_09238__699 VPWR VGND net699 sg13g2_tiehi
XFILLER_42_897 VPWR VGND sg13g2_fill_1
XFILLER_96_514 VPWR VGND sg13g2_decap_4
XFILLER_2_971 VPWR VGND sg13g2_decap_8
XFILLER_39_6 VPWR VGND sg13g2_fill_1
Xinput7 ui_in[5] net7 VPWR VGND sg13g2_buf_1
XFILLER_64_400 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_4_clk_regs clknet_5_2__leaf_clk_regs clknet_leaf_4_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_37_625 VPWR VGND sg13g2_decap_8
X_08117__577 VPWR VGND net577 sg13g2_tiehi
X_05610_ VGND VPWR net1067 _02277_ _00028_ _02278_ sg13g2_a21oi_1
X_06590_ net3504 net1154 _02650_ VPWR VGND sg13g2_nor2_1
XFILLER_33_820 VPWR VGND sg13g2_fill_1
X_05541_ _02227_ net3643 net1070 VPWR VGND sg13g2_nand2_1
X_08260_ net417 VGND VPWR _00341_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[27\]
+ clknet_leaf_58_clk_regs sg13g2_dfrbpq_1
X_05472_ i_exotiny._1611_\[3\] net1281 net3702 net13 VPWR VGND sg13g2_and3_1
X_08191_ net486 VGND VPWR _00272_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[22\]
+ clknet_leaf_68_clk_regs sg13g2_dfrbpq_1
X_07211_ net1905 net1088 _02967_ VPWR VGND sg13g2_nor2_1
X_07142_ VGND VPWR net1159 _02948_ _02947_ net1142 sg13g2_a21oi_2
XFILLER_106_608 VPWR VGND sg13g2_decap_8
X_07073_ i_exotiny._0015_\[1\] net3368 net916 _00828_ VPWR VGND sg13g2_mux2_1
X_06024_ VGND VPWR i_exotiny._1615_\[3\] net1103 _00214_ _02506_ sg13g2_a21oi_1
XFILLER_102_825 VPWR VGND sg13g2_decap_8
XFILLER_99_374 VPWR VGND sg13g2_decap_8
XFILLER_101_324 VPWR VGND sg13g2_decap_8
X_07975_ net116 VGND VPWR i_exotiny._1611_\[3\] i_exotiny._0369_\[27\] clknet_leaf_11_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_74_219 VPWR VGND sg13g2_fill_2
X_06926_ net2408 net2783 net925 _00705_ VPWR VGND sg13g2_mux2_1
X_06857_ net1872 net1189 _02868_ VPWR VGND sg13g2_nor2_1
X_05808_ net2484 i_exotiny._0018_\[0\] net1056 _00080_ VPWR VGND sg13g2_mux2_1
X_06788_ VGND VPWR net1098 _02809_ _00674_ _02810_ sg13g2_a21oi_1
X_09055__927 VPWR VGND net1347 sg13g2_tiehi
X_05739_ i_exotiny.i_wb_spi.cnt_hbit_r\[5\] _02368_ _02376_ VPWR VGND sg13g2_nor2_1
X_08527_ net153 VGND VPWR net2225 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[15\]
+ clknet_leaf_182_clk_regs sg13g2_dfrbpq_1
X_08458_ net222 VGND VPWR net2551 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[10\]
+ clknet_leaf_114_clk_regs sg13g2_dfrbpq_1
X_07409_ VGND VPWR i_exotiny._0369_\[14\] _03050_ _03059_ _03052_ sg13g2_a21oi_1
XFILLER_13_1025 VPWR VGND sg13g2_decap_4
X_08389_ net289 VGND VPWR _00470_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[27\]
+ clknet_leaf_140_clk_regs sg13g2_dfrbpq_1
Xclkbuf_leaf_74_clk_regs clknet_5_26__leaf_clk_regs clknet_leaf_74_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_3_746 VPWR VGND sg13g2_decap_8
XFILLER_105_685 VPWR VGND sg13g2_decap_8
XFILLER_104_173 VPWR VGND sg13g2_decap_8
XFILLER_66_709 VPWR VGND sg13g2_fill_2
X_09240__567 VPWR VGND net567 sg13g2_tiehi
XFILLER_76_98 VPWR VGND sg13g2_fill_2
XFILLER_19_669 VPWR VGND sg13g2_fill_1
XFILLER_61_425 VPWR VGND sg13g2_fill_1
X_08690__1298 VPWR VGND net1718 sg13g2_tiehi
XFILLER_18_179 VPWR VGND sg13g2_fill_1
XFILLER_15_864 VPWR VGND sg13g2_fill_2
Xclkbuf_4_4_0_clk_regs clknet_0_clk_regs clknet_4_4_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_97_856 VPWR VGND sg13g2_decap_8
XFILLER_96_322 VPWR VGND sg13g2_decap_8
Xhold1708 i_exotiny._1160_\[21\] VPWR VGND net3535 sg13g2_dlygate4sd3_1
X_07760_ net3170 net2404 net991 _01245_ VPWR VGND sg13g2_mux2_1
Xhold1719 _01083_ VPWR VGND net3546 sg13g2_dlygate4sd3_1
XFILLER_37_400 VPWR VGND sg13g2_fill_2
X_04972_ _01704_ i_exotiny._0315_\[5\] _01703_ VPWR VGND sg13g2_xnor2_1
XFILLER_96_399 VPWR VGND sg13g2_fill_2
XFILLER_77_580 VPWR VGND sg13g2_fill_2
X_06711_ _01390_ net1233 i_exotiny._0315_\[4\] _02745_ VGND VPWR _02721_ sg13g2_nor4_2
XFILLER_49_293 VPWR VGND sg13g2_fill_2
X_07691_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[26\]
+ net2172 net1000 _01193_ VPWR VGND sg13g2_mux2_1
X_06642_ net1198 _02683_ _02684_ _00654_ VPWR VGND sg13g2_nor3_1
X_06573_ net1200 _02637_ _02638_ _00631_ VPWR VGND sg13g2_nor3_1
X_08312_ net366 VGND VPWR net3286 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[14\]
+ clknet_leaf_76_clk_regs sg13g2_dfrbpq_1
XFILLER_80_789 VPWR VGND sg13g2_fill_1
X_09292_ net1815 VGND VPWR net2260 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[18\]
+ clknet_leaf_171_clk_regs sg13g2_dfrbpq_1
X_05524_ net1276 i_exotiny._0315_\[14\] _02213_ VPWR VGND sg13g2_nor2b_1
X_08243_ net434 VGND VPWR _00324_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[10\]
+ clknet_leaf_48_clk_regs sg13g2_dfrbpq_1
X_05455_ VPWR VGND i_exotiny._1618_\[2\] _02161_ _02140_ i_exotiny._1614_\[2\] _02162_
+ _02135_ sg13g2_a221oi_1
X_05386_ VPWR i_exotiny._2055_\[2\] net3327 VGND sg13g2_inv_1
X_08174_ net503 VGND VPWR _00255_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[5\]
+ clknet_leaf_112_clk_regs sg13g2_dfrbpq_1
X_04658__1 VPWR net1827 clknet_1_0__leaf_clk VGND sg13g2_inv_1
XFILLER_106_405 VPWR VGND sg13g2_decap_8
X_07125_ net1287 net1867 _00875_ VPWR VGND sg13g2_and2_1
X_07056_ net3275 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[22\]
+ net1017 _00817_ VPWR VGND sg13g2_mux2_1
X_08198__479 VPWR VGND net479 sg13g2_tiehi
X_08888__1094 VPWR VGND net1514 sg13g2_tiehi
X_06007_ net2156 _02497_ net1048 _00206_ VPWR VGND sg13g2_mux2_1
XFILLER_0_749 VPWR VGND sg13g2_decap_8
XFILLER_87_388 VPWR VGND sg13g2_fill_1
XFILLER_75_517 VPWR VGND sg13g2_decap_4
XFILLER_29_901 VPWR VGND sg13g2_fill_2
XFILLER_101_198 VPWR VGND sg13g2_decap_8
X_07958_ net698 VGND VPWR net1993 i_exotiny.i_wb_spi.cnt_hbit_r\[3\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_68_591 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_121_clk_regs clknet_5_22__leaf_clk_regs clknet_leaf_121_clk_regs VPWR
+ VGND sg13g2_buf_8
X_06909_ _02909_ i_exotiny._1586_ i_exotiny.i_rstctl.cnt\[3\] VPWR VGND sg13g2_nand2_1
X_07889_ net2190 net2779 net980 _01356_ VPWR VGND sg13g2_mux2_1
XFILLER_15_149 VPWR VGND sg13g2_fill_2
XFILLER_43_447 VPWR VGND sg13g2_fill_1
XFILLER_62_45 VPWR VGND sg13g2_fill_1
XFILLER_12_845 VPWR VGND sg13g2_fill_2
X_08675__1313 VPWR VGND net1733 sg13g2_tiehi
X_08107__587 VPWR VGND net587 sg13g2_tiehi
XFILLER_106_972 VPWR VGND sg13g2_decap_8
XFILLER_87_31 VPWR VGND sg13g2_fill_2
XFILLER_78_300 VPWR VGND sg13g2_fill_1
XFILLER_93_303 VPWR VGND sg13g2_decap_8
XFILLER_93_325 VPWR VGND sg13g2_decap_8
XFILLER_4_1023 VPWR VGND sg13g2_decap_4
XFILLER_62_701 VPWR VGND sg13g2_fill_1
XFILLER_35_904 VPWR VGND sg13g2_fill_2
XFILLER_59_1025 VPWR VGND sg13g2_decap_4
X_09038__944 VPWR VGND net1364 sg13g2_tiehi
XFILLER_99_5 VPWR VGND sg13g2_fill_2
Xinput10 uio_in[0] net10 VPWR VGND sg13g2_buf_2
X_05240_ _01612_ _01966_ _01967_ _01968_ VPWR VGND sg13g2_nor3_1
X_05171_ _01825_ _01898_ _01899_ _01900_ VPWR VGND sg13g2_or3_1
Xhold827 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[5\]
+ VPWR VGND net2654 sg13g2_dlygate4sd3_1
Xhold816 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[17\]
+ VPWR VGND net2643 sg13g2_dlygate4sd3_1
X_09298__1347 VPWR VGND net1767 sg13g2_tiehi
Xhold805 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[11\]
+ VPWR VGND net2632 sg13g2_dlygate4sd3_1
XFILLER_104_909 VPWR VGND sg13g2_decap_8
Xhold849 _00144_ VPWR VGND net2676 sg13g2_dlygate4sd3_1
Xhold838 _00312_ VPWR VGND net2665 sg13g2_dlygate4sd3_1
X_08930_ net1472 VGND VPWR net3072 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[28\]
+ clknet_leaf_65_clk_regs sg13g2_dfrbpq_1
X_08861_ net1545 VGND VPWR net3534 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[28\]
+ clknet_leaf_184_clk_regs sg13g2_dfrbpq_1
XFILLER_35_0 VPWR VGND sg13g2_decap_4
Xhold1516 i_exotiny._0035_\[2\] VPWR VGND net3343 sg13g2_dlygate4sd3_1
Xhold1505 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[22\]
+ VPWR VGND net3332 sg13g2_dlygate4sd3_1
X_07812_ net2733 net2704 net891 _01291_ VPWR VGND sg13g2_mux2_1
Xhold1527 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[13\]
+ VPWR VGND net3354 sg13g2_dlygate4sd3_1
Xhold1549 _01294_ VPWR VGND net3376 sg13g2_dlygate4sd3_1
Xhold1538 _00837_ VPWR VGND net3365 sg13g2_dlygate4sd3_1
X_08792_ net1616 VGND VPWR _00850_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[23\]
+ clknet_leaf_164_clk_regs sg13g2_dfrbpq_1
X_07743_ _01231_ _03205_ _03208_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_230 VPWR VGND sg13g2_fill_2
X_04955_ _01532_ i_exotiny._0315_\[7\] net1201 _01687_ VPWR VGND sg13g2_mux2_1
X_08753__1235 VPWR VGND net1655 sg13g2_tiehi
XFILLER_53_723 VPWR VGND sg13g2_fill_2
X_07674_ net2301 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[13\]
+ net998 _01176_ VPWR VGND sg13g2_mux2_1
X_04886_ net1222 _01616_ _01617_ _01618_ VPWR VGND sg13g2_nor3_2
XFILLER_52_233 VPWR VGND sg13g2_fill_2
X_06625_ i_exotiny._0314_\[21\] net1159 _02673_ VPWR VGND sg13g2_nor2_1
X_06556_ net1261 net3596 net1216 _00623_ VPWR VGND sg13g2_mux2_1
X_06487_ net3021 net3298 net1026 _00568_ VPWR VGND sg13g2_mux2_1
X_09275_ net71 VGND VPWR net2372 i_exotiny._0021_\[1\] clknet_leaf_178_clk_regs sg13g2_dfrbpq_2
XFILLER_20_141 VPWR VGND sg13g2_fill_2
XFILLER_21_664 VPWR VGND sg13g2_fill_1
X_05507_ _02200_ net2125 net1069 VPWR VGND sg13g2_nand2_1
XFILLER_32_37 VPWR VGND sg13g2_decap_8
X_05438_ _02147_ _02146_ i_exotiny._1616_\[0\] _02145_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data[0]
+ VPWR VGND sg13g2_a22oi_1
X_08226_ net451 VGND VPWR net2390 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[25\]
+ clknet_leaf_153_clk_regs sg13g2_dfrbpq_1
XFILLER_32_48 VPWR VGND sg13g2_fill_1
X_08157_ net521 VGND VPWR net2392 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[21\]
+ clknet_leaf_133_clk_regs sg13g2_dfrbpq_1
XFILLER_106_202 VPWR VGND sg13g2_decap_8
X_05369_ _02078_ _02088_ _02089_ _02090_ _02091_ VPWR VGND sg13g2_nor4_1
X_07108_ _02381_ net1111 net1227 _02946_ VPWR VGND sg13g2_a21o_1
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
X_08975__1007 VPWR VGND net1427 sg13g2_tiehi
X_08088_ net606 VGND VPWR _00169_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[25\]
+ clknet_leaf_92_clk_regs sg13g2_dfrbpq_1
XFILLER_106_279 VPWR VGND sg13g2_decap_8
X_07039_ net2293 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[5\]
+ net1015 _00800_ VPWR VGND sg13g2_mux2_1
XFILLER_103_986 VPWR VGND sg13g2_decap_8
XFILLER_102_441 VPWR VGND sg13g2_decap_8
XFILLER_87_130 VPWR VGND sg13g2_fill_1
XFILLER_28_285 VPWR VGND sg13g2_fill_1
X_08624__1352 VPWR VGND net1772 sg13g2_tiehi
XFILLER_4_841 VPWR VGND sg13g2_decap_8
X_08831__1157 VPWR VGND net1577 sg13g2_tiehi
XFILLER_98_439 VPWR VGND sg13g2_decap_8
XFILLER_78_152 VPWR VGND sg13g2_fill_1
Xfanout1130 net1131 net1130 VPWR VGND sg13g2_buf_8
Xfanout1141 net1142 net1141 VPWR VGND sg13g2_buf_8
Xfanout1152 net1153 net1152 VPWR VGND sg13g2_buf_8
Xfanout1163 net1164 net1163 VPWR VGND sg13g2_buf_8
Xfanout1174 _01435_ net1174 VPWR VGND sg13g2_buf_8
XFILLER_66_347 VPWR VGND sg13g2_fill_1
Xfanout1185 net1187 net1185 VPWR VGND sg13g2_buf_8
Xfanout1196 net1197 net1196 VPWR VGND sg13g2_buf_8
X_04740_ VGND VPWR i_exotiny._1306_ _01476_ _01495_ net1893 sg13g2_a21oi_1
XFILLER_47_561 VPWR VGND sg13g2_fill_2
XFILLER_19_296 VPWR VGND sg13g2_fill_1
X_08188__489 VPWR VGND net489 sg13g2_tiehi
XFILLER_62_553 VPWR VGND sg13g2_fill_2
XFILLER_34_255 VPWR VGND sg13g2_fill_1
XFILLER_35_767 VPWR VGND sg13g2_fill_1
X_04671_ net1248 net1254 _01432_ VPWR VGND sg13g2_nor2_1
X_06410_ _02590_ VPWR _00514_ VGND _02219_ _02592_ sg13g2_o21ai_1
XFILLER_97_2 VPWR VGND sg13g2_fill_1
XFILLER_34_277 VPWR VGND sg13g2_fill_1
X_07390_ net1955 net1077 _03043_ VPWR VGND sg13g2_nor2_1
X_06341_ _02563_ net2971 net1033 _00474_ VPWR VGND sg13g2_mux2_1
X_09060_ net1342 VGND VPWR net1831 i_exotiny.i_wdg_top.clk_div_inst.cnt\[0\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
X_06272_ net2402 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[4\]
+ net942 _00415_ VPWR VGND sg13g2_mux2_1
X_08011_ net684 VGND VPWR net2153 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[12\]
+ clknet_leaf_62_clk_regs sg13g2_dfrbpq_1
X_05223_ _01951_ _01627_ i_exotiny._0028_\[1\] _01622_ i_exotiny._0023_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold602 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[24\]
+ VPWR VGND net2429 sg13g2_dlygate4sd3_1
XFILLER_104_706 VPWR VGND sg13g2_decap_8
Xhold635 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[6\]
+ VPWR VGND net2462 sg13g2_dlygate4sd3_1
Xhold624 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[6\]
+ VPWR VGND net2451 sg13g2_dlygate4sd3_1
Xhold613 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[11\]
+ VPWR VGND net2440 sg13g2_dlygate4sd3_1
X_05154_ _01643_ VPWR _01884_ VGND net1255 i_exotiny._0018_\[2\] sg13g2_o21ai_1
X_08807__1181 VPWR VGND net1601 sg13g2_tiehi
Xhold668 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[31\]
+ VPWR VGND net2495 sg13g2_dlygate4sd3_1
Xhold679 _00175_ VPWR VGND net2506 sg13g2_dlygate4sd3_1
Xhold646 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[21\]
+ VPWR VGND net2473 sg13g2_dlygate4sd3_1
Xhold657 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[4\]
+ VPWR VGND net2484 sg13g2_dlygate4sd3_1
X_05085_ _01816_ _01467_ _01430_ VPWR VGND sg13g2_nand2b_1
XFILLER_103_227 VPWR VGND sg13g2_decap_8
XFILLER_98_951 VPWR VGND sg13g2_decap_8
X_08913_ net1489 VGND VPWR _00971_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[11\]
+ clknet_leaf_66_clk_regs sg13g2_dfrbpq_1
Xhold2003 i_exotiny._1757_ VPWR VGND net3830 sg13g2_dlygate4sd3_1
XFILLER_97_450 VPWR VGND sg13g2_fill_2
Xhold2014 i_exotiny._3871_ VPWR VGND net3841 sg13g2_dlygate4sd3_1
XFILLER_100_945 VPWR VGND sg13g2_decap_8
Xhold1302 i_exotiny._0017_\[1\] VPWR VGND net3129 sg13g2_dlygate4sd3_1
Xhold1324 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[24\]
+ VPWR VGND net3151 sg13g2_dlygate4sd3_1
X_08844_ net1562 VGND VPWR _00902_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[11\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
Xhold1313 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[7\]
+ VPWR VGND net3140 sg13g2_dlygate4sd3_1
Xhold1335 _00344_ VPWR VGND net3162 sg13g2_dlygate4sd3_1
Xhold1368 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[15\]
+ VPWR VGND net3195 sg13g2_dlygate4sd3_1
Xhold1346 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[31\]
+ VPWR VGND net3173 sg13g2_dlygate4sd3_1
X_05987_ net2595 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[17\]
+ net1050 _00189_ VPWR VGND sg13g2_mux2_1
X_08775_ net1633 VGND VPWR net3074 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[6\]
+ clknet_leaf_158_clk_regs sg13g2_dfrbpq_1
Xhold1357 _00786_ VPWR VGND net3184 sg13g2_dlygate4sd3_1
Xhold1379 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[30\]
+ VPWR VGND net3206 sg13g2_dlygate4sd3_1
X_07726_ net2387 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[23\]
+ net993 _01222_ VPWR VGND sg13g2_mux2_1
XFILLER_27_59 VPWR VGND sg13g2_fill_2
X_04938_ _01668_ _01669_ _01667_ _01670_ VPWR VGND sg13g2_nand3_1
X_07657_ net3006 net882 _03187_ _03190_ VPWR VGND sg13g2_mux2_1
X_04869_ net1271 net1267 net1268 _01601_ VPWR VGND sg13g2_nor3_2
X_07588_ net1204 net1914 _03163_ _01121_ VPWR VGND sg13g2_nor3_1
X_06608_ net3243 net1155 _02662_ VPWR VGND sg13g2_nor2_1
X_06539_ net3031 net886 _02620_ _02622_ VPWR VGND sg13g2_mux2_1
XFILLER_43_58 VPWR VGND sg13g2_fill_1
X_09258_ net509 VGND VPWR _01313_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[16\]
+ clknet_leaf_128_clk_regs sg13g2_dfrbpq_1
X_09189_ net792 VGND VPWR net2744 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[11\]
+ clknet_leaf_77_clk_regs sg13g2_dfrbpq_1
XFILLER_5_638 VPWR VGND sg13g2_fill_1
X_08209_ net468 VGND VPWR net2763 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[8\]
+ clknet_leaf_150_clk_regs sg13g2_dfrbpq_1
X_08004__691 VPWR VGND net691 sg13g2_tiehi
XFILLER_1_866 VPWR VGND sg13g2_decap_8
X_09028__954 VPWR VGND net1374 sg13g2_tiehi
XFILLER_103_783 VPWR VGND sg13g2_decap_8
XFILLER_89_995 VPWR VGND sg13g2_decap_8
XFILLER_48_347 VPWR VGND sg13g2_fill_2
Xhold1880 i_exotiny._1711_ VPWR VGND net3707 sg13g2_dlygate4sd3_1
Xhold1891 _00680_ VPWR VGND net3718 sg13g2_dlygate4sd3_1
XFILLER_29_594 VPWR VGND sg13g2_fill_1
XFILLER_32_737 VPWR VGND sg13g2_fill_1
X_08011__684 VPWR VGND net684 sg13g2_tiehi
XFILLER_13_962 VPWR VGND sg13g2_decap_8
X_09035__947 VPWR VGND net1367 sg13g2_tiehi
XFILLER_9_988 VPWR VGND sg13g2_decap_8
X_09081__901 VPWR VGND net1321 sg13g2_tiehi
X_05910_ net2903 net2975 net973 _00127_ VPWR VGND sg13g2_mux2_1
X_06890_ VGND VPWR i_exotiny._1618_\[3\] net1128 _02896_ _02895_ sg13g2_a21oi_1
XFILLER_95_954 VPWR VGND sg13g2_decap_8
X_05841_ _02430_ _01497_ _02048_ VPWR VGND sg13g2_nand2_1
XFILLER_54_317 VPWR VGND sg13g2_fill_2
X_05772_ _02399_ net1126 _01377_ net1144 net3785 VPWR VGND sg13g2_a22oi_1
X_08560_ net84 VGND VPWR net3383 i_exotiny._0314_\[5\] clknet_leaf_5_clk_regs sg13g2_dfrbpq_2
XFILLER_63_884 VPWR VGND sg13g2_fill_2
X_08491_ net189 VGND VPWR _00565_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[11\]
+ clknet_leaf_106_clk_regs sg13g2_dfrbpq_1
X_07511_ net2099 net2841 net901 _01094_ VPWR VGND sg13g2_mux2_1
XFILLER_23_715 VPWR VGND sg13g2_fill_2
X_04723_ VGND VPWR _01455_ _01480_ _00004_ net1197 sg13g2_a21oi_1
X_04654_ VPWR _01416_ net1951 VGND sg13g2_inv_1
XFILLER_22_203 VPWR VGND sg13g2_fill_1
X_07442_ _03084_ net1149 _03083_ net1209 i_exotiny._1160_\[22\] VPWR VGND sg13g2_a22oi_1
X_07373_ VGND VPWR net1078 _03029_ _01039_ _03030_ sg13g2_a21oi_1
X_06324_ net2949 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[18\]
+ net1035 _00461_ VPWR VGND sg13g2_mux2_1
X_09112_ net870 VGND VPWR net2183 i_exotiny._0030_\[0\] clknet_leaf_157_clk_regs sg13g2_dfrbpq_2
XFILLER_30_280 VPWR VGND sg13g2_fill_1
X_09267__93 VPWR VGND net93 sg13g2_tiehi
X_06255_ net3164 net3409 net1039 _00404_ VPWR VGND sg13g2_mux2_1
X_09043_ net1570 VGND VPWR net2025 i_exotiny._0315_\[31\] clknet_leaf_2_clk_regs sg13g2_dfrbpq_2
X_06186_ _02472_ net3212 _02533_ _02538_ VPWR VGND sg13g2_mux2_1
Xhold410 _01155_ VPWR VGND net2237 sg13g2_dlygate4sd3_1
X_05206_ _01930_ _01933_ _01934_ VPWR VGND sg13g2_nor2_1
Xhold443 _00482_ VPWR VGND net2270 sg13g2_dlygate4sd3_1
Xhold421 _00094_ VPWR VGND net2248 sg13g2_dlygate4sd3_1
Xhold454 _00746_ VPWR VGND net2281 sg13g2_dlygate4sd3_1
Xhold432 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[22\]
+ VPWR VGND net2259 sg13g2_dlygate4sd3_1
X_05137_ _01849_ _01861_ _01755_ _01867_ VPWR VGND _01866_ sg13g2_nand4_1
Xhold487 _00821_ VPWR VGND net2314 sg13g2_dlygate4sd3_1
Xhold465 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[18\]
+ VPWR VGND net2292 sg13g2_dlygate4sd3_1
Xhold476 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[7\]
+ VPWR VGND net2303 sg13g2_dlygate4sd3_1
Xfanout912 _02979_ net912 VPWR VGND sg13g2_buf_8
Xhold498 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[12\]
+ VPWR VGND net2325 sg13g2_dlygate4sd3_1
Xfanout901 net902 net901 VPWR VGND sg13g2_buf_8
Xfanout934 net936 net934 VPWR VGND sg13g2_buf_8
X_05068_ _01800_ _01789_ i_exotiny._0024_\[3\] _01765_ i_exotiny._0027_\[3\] VPWR
+ VGND sg13g2_a22oi_1
Xfanout923 _02929_ net923 VPWR VGND sg13g2_buf_2
Xfanout967 net971 net967 VPWR VGND sg13g2_buf_8
Xfanout956 net957 net956 VPWR VGND sg13g2_buf_8
Xfanout945 net949 net945 VPWR VGND sg13g2_buf_8
X_08827_ net1581 VGND VPWR _00885_ i_exotiny.i_wb_spi.state_r\[26\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
Xfanout989 _03211_ net989 VPWR VGND sg13g2_buf_1
XFILLER_86_976 VPWR VGND sg13g2_decap_8
Xhold1121 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[24\]
+ VPWR VGND net2948 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_99_clk_regs clknet_5_29__leaf_clk_regs clknet_leaf_99_clk_regs VPWR VGND
+ sg13g2_buf_8
Xfanout978 net980 net978 VPWR VGND sg13g2_buf_8
Xhold1132 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[5\]
+ VPWR VGND net2959 sg13g2_dlygate4sd3_1
Xhold1110 _00856_ VPWR VGND net2937 sg13g2_dlygate4sd3_1
Xhold1143 _00154_ VPWR VGND net2970 sg13g2_dlygate4sd3_1
XFILLER_79_1028 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_28_clk_regs clknet_5_9__leaf_clk_regs clknet_leaf_28_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold1176 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[12\]
+ VPWR VGND net3003 sg13g2_dlygate4sd3_1
Xhold1165 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[4\]
+ VPWR VGND net2992 sg13g2_dlygate4sd3_1
Xhold1154 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[21\]
+ VPWR VGND net2981 sg13g2_dlygate4sd3_1
X_08758_ net1650 VGND VPWR net2574 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[21\]
+ clknet_leaf_87_clk_regs sg13g2_dfrbpq_1
Xhold1187 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[16\]
+ VPWR VGND net3014 sg13g2_dlygate4sd3_1
Xhold1198 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[18\]
+ VPWR VGND net3025 sg13g2_dlygate4sd3_1
X_08689_ net1719 VGND VPWR _00747_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[16\]
+ clknet_leaf_102_clk_regs sg13g2_dfrbpq_1
X_07709_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[10\]
+ net2724 net996 _01205_ VPWR VGND sg13g2_mux2_1
XFILLER_14_737 VPWR VGND sg13g2_fill_1
XFILLER_10_998 VPWR VGND sg13g2_decap_8
XFILLER_6_969 VPWR VGND sg13g2_decap_8
X_08178__499 VPWR VGND net499 sg13g2_tiehi
XFILLER_88_291 VPWR VGND sg13g2_fill_2
XFILLER_37_807 VPWR VGND sg13g2_decap_4
XFILLER_92_935 VPWR VGND sg13g2_decap_8
XFILLER_36_306 VPWR VGND sg13g2_fill_1
XFILLER_36_339 VPWR VGND sg13g2_fill_1
XFILLER_17_586 VPWR VGND sg13g2_decap_4
XFILLER_32_523 VPWR VGND sg13g2_fill_1
XFILLER_32_534 VPWR VGND sg13g2_decap_4
X_08970__1012 VPWR VGND net1432 sg13g2_tiehi
XFILLER_81_5 VPWR VGND sg13g2_fill_1
X_06040_ net2240 net2464 net964 _00225_ VPWR VGND sg13g2_mux2_1
XFILLER_5_980 VPWR VGND sg13g2_decap_8
XFILLER_101_506 VPWR VGND sg13g2_decap_8
X_08688__1300 VPWR VGND net1720 sg13g2_tiehi
X_07991_ net132 VGND VPWR net3750 i_exotiny._0369_\[1\] clknet_leaf_11_clk_regs sg13g2_dfrbpq_1
X_06942_ net2278 net3056 net925 _00721_ VPWR VGND sg13g2_mux2_1
XFILLER_95_784 VPWR VGND sg13g2_fill_1
X_06873_ net3668 net1094 _02882_ VPWR VGND sg13g2_nor2_1
X_05824_ net2453 net2152 net1053 _00096_ VPWR VGND sg13g2_mux2_1
X_08612_ net1784 VGND VPWR net3502 i_exotiny._1616_\[0\] clknet_leaf_22_clk_regs sg13g2_dfrbpq_2
X_05755_ _02388_ _02385_ net3399 VPWR VGND sg13g2_nand2b_1
X_08543_ net113 VGND VPWR net2492 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[31\]
+ clknet_leaf_182_clk_regs sg13g2_dfrbpq_1
XFILLER_36_873 VPWR VGND sg13g2_fill_2
XFILLER_82_489 VPWR VGND sg13g2_fill_1
XFILLER_23_501 VPWR VGND sg13g2_fill_1
XFILLER_23_512 VPWR VGND sg13g2_fill_2
X_04706_ _01464_ net1249 _01462_ _01463_ VPWR VGND sg13g2_and3_2
X_05686_ VGND VPWR net1063 _02335_ _00047_ _02333_ sg13g2_a21oi_1
X_08474_ net206 VGND VPWR _00548_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[26\]
+ clknet_leaf_114_clk_regs sg13g2_dfrbpq_1
XFILLER_51_854 VPWR VGND sg13g2_fill_2
XFILLER_24_38 VPWR VGND sg13g2_fill_1
X_04637_ VPWR _01399_ i_exotiny._2034_\[1\] VGND sg13g2_inv_1
X_09018__964 VPWR VGND net1384 sg13g2_tiehi
X_07425_ VGND VPWR i_exotiny._0369_\[18\] net1147 _03071_ _03052_ sg13g2_a21oi_1
Xclkbuf_leaf_146_clk_regs clknet_5_16__leaf_clk_regs clknet_leaf_146_clk_regs VPWR
+ VGND sg13g2_buf_8
X_07356_ VGND VPWR net1078 _03017_ _01035_ _03012_ sg13g2_a21oi_1
X_07287_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[12\]
+ net2715 net910 _01004_ VPWR VGND sg13g2_mux2_1
X_06307_ net2465 i_exotiny._0014_\[1\] net1033 _00444_ VPWR VGND sg13g2_mux2_1
XFILLER_40_26 VPWR VGND sg13g2_fill_1
X_06238_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[12\]
+ net2986 net1040 _00387_ VPWR VGND sg13g2_mux2_1
X_09026_ net1376 VGND VPWR net3548 i_exotiny._0315_\[14\] clknet_leaf_167_clk_regs
+ sg13g2_dfrbpq_1
X_08394__534 VPWR VGND net534 sg13g2_tiehi
XFILLER_3_928 VPWR VGND sg13g2_decap_8
Xhold240 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[13\]
+ VPWR VGND net2067 sg13g2_dlygate4sd3_1
X_06169_ net2873 net3096 net951 _00331_ VPWR VGND sg13g2_mux2_1
Xhold251 _01049_ VPWR VGND net2078 sg13g2_dlygate4sd3_1
Xhold262 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[9\]
+ VPWR VGND net2089 sg13g2_dlygate4sd3_1
XFILLER_105_867 VPWR VGND sg13g2_decap_8
XFILLER_104_355 VPWR VGND sg13g2_decap_8
Xhold284 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[26\]
+ VPWR VGND net2111 sg13g2_dlygate4sd3_1
Xhold273 _01098_ VPWR VGND net2100 sg13g2_dlygate4sd3_1
Xhold295 _01323_ VPWR VGND net2122 sg13g2_dlygate4sd3_1
X_08001__694 VPWR VGND net694 sg13g2_tiehi
X_08848__1138 VPWR VGND net1558 sg13g2_tiehi
XFILLER_105_30 VPWR VGND sg13g2_decap_4
X_09025__957 VPWR VGND net1377 sg13g2_tiehi
XFILLER_46_615 VPWR VGND sg13g2_fill_1
XFILLER_45_136 VPWR VGND sg13g2_fill_1
XFILLER_42_821 VPWR VGND sg13g2_fill_1
X_09071__911 VPWR VGND net1331 sg13g2_tiehi
X_08766__1222 VPWR VGND net1642 sg13g2_tiehi
XFILLER_5_243 VPWR VGND sg13g2_fill_1
X_08799__1189 VPWR VGND net1609 sg13g2_tiehi
XFILLER_2_950 VPWR VGND sg13g2_decap_8
XFILLER_7_1010 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[6] net8 VPWR VGND sg13g2_buf_1
XFILLER_91_231 VPWR VGND sg13g2_fill_2
XFILLER_91_297 VPWR VGND sg13g2_fill_1
X_05540_ _02218_ VPWR i_exotiny._1611_\[25\] VGND _02219_ _02225_ sg13g2_o21ai_1
XFILLER_45_692 VPWR VGND sg13g2_decap_8
X_05471_ net1076 VPWR i_exotiny._1611_\[2\] VGND _01405_ _01543_ sg13g2_o21ai_1
X_07210_ VGND VPWR _01414_ net1089 _00940_ _02966_ sg13g2_a21oi_1
X_08190_ net487 VGND VPWR net2594 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[21\]
+ clknet_leaf_111_clk_regs sg13g2_dfrbpq_1
X_07141_ _02419_ _02532_ _02947_ VPWR VGND sg13g2_nor2_2
X_07072_ net3063 net3000 net914 _00827_ VPWR VGND sg13g2_mux2_1
X_06023_ net3543 net1103 _02506_ VPWR VGND sg13g2_nor2_1
XFILLER_102_804 VPWR VGND sg13g2_decap_8
XFILLER_99_353 VPWR VGND sg13g2_decap_8
XFILLER_101_303 VPWR VGND sg13g2_decap_8
XFILLER_87_504 VPWR VGND sg13g2_decap_4
X_07974_ net115 VGND VPWR i_exotiny._1611_\[2\] i_exotiny._0369_\[26\] clknet_leaf_21_clk_regs
+ sg13g2_dfrbpq_1
X_09292__1395 VPWR VGND net1815 sg13g2_tiehi
X_06925_ net2524 net2856 net924 _00704_ VPWR VGND sg13g2_mux2_1
XFILLER_67_283 VPWR VGND sg13g2_fill_1
X_06856_ VGND VPWR net1094 _02866_ _00685_ _02867_ sg13g2_a21oi_1
XFILLER_55_434 VPWR VGND sg13g2_decap_8
XFILLER_28_626 VPWR VGND sg13g2_fill_2
XFILLER_71_905 VPWR VGND sg13g2_fill_2
XFILLER_55_456 VPWR VGND sg13g2_decap_4
X_05807_ VGND VPWR _02414_ _02424_ net1142 _02421_ sg13g2_a21oi_2
X_06787_ net3622 net1098 _02810_ VPWR VGND sg13g2_nor2_1
XFILLER_42_106 VPWR VGND sg13g2_fill_1
X_05738_ _02373_ VPWR _02375_ VGND i_exotiny.i_wb_regs.spi_size_o\[0\] i_exotiny.i_wb_regs.spi_size_o\[1\]
+ sg13g2_o21ai_1
X_08526_ net154 VGND VPWR net2185 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[14\]
+ clknet_leaf_183_clk_regs sg13g2_dfrbpq_1
XFILLER_23_331 VPWR VGND sg13g2_fill_1
X_05669_ VGND VPWR i_exotiny._1617_\[1\] net1122 _02323_ _02322_ sg13g2_a21oi_1
XFILLER_24_887 VPWR VGND sg13g2_fill_2
X_08457_ net223 VGND VPWR net2233 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[9\]
+ clknet_leaf_158_clk_regs sg13g2_dfrbpq_1
XFILLER_11_548 VPWR VGND sg13g2_fill_2
X_07408_ net2040 net1215 _03058_ VPWR VGND sg13g2_nor2_1
XFILLER_7_519 VPWR VGND sg13g2_fill_1
XFILLER_13_1004 VPWR VGND sg13g2_decap_8
X_08388_ net290 VGND VPWR _00469_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[26\]
+ clknet_leaf_140_clk_regs sg13g2_dfrbpq_1
X_07339_ _03002_ VPWR _03003_ VGND i_exotiny._0369_\[7\] _02995_ sg13g2_o21ai_1
X_09009_ net1393 VGND VPWR _01067_ i_exotiny._0079_\[2\] clknet_leaf_159_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_105_664 VPWR VGND sg13g2_decap_8
XFILLER_2_224 VPWR VGND sg13g2_fill_2
X_09262__237 VPWR VGND net237 sg13g2_tiehi
XFILLER_104_152 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_43_clk_regs clknet_5_10__leaf_clk_regs clknet_leaf_43_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_78_504 VPWR VGND sg13g2_fill_1
XFILLER_59_751 VPWR VGND sg13g2_fill_1
XFILLER_101_892 VPWR VGND sg13g2_decap_8
XFILLER_46_434 VPWR VGND sg13g2_fill_1
XFILLER_74_776 VPWR VGND sg13g2_fill_1
XFILLER_18_147 VPWR VGND sg13g2_fill_1
XFILLER_33_117 VPWR VGND sg13g2_fill_2
XFILLER_92_98 VPWR VGND sg13g2_fill_2
XFILLER_10_581 VPWR VGND sg13g2_fill_1
XFILLER_6_552 VPWR VGND sg13g2_fill_2
X_08123__571 VPWR VGND net571 sg13g2_tiehi
XFILLER_97_835 VPWR VGND sg13g2_decap_8
XFILLER_96_301 VPWR VGND sg13g2_decap_8
XFILLER_69_515 VPWR VGND sg13g2_fill_1
XFILLER_37_4 VPWR VGND sg13g2_decap_8
XFILLER_96_378 VPWR VGND sg13g2_decap_8
X_04971_ _01420_ _01423_ i_exotiny._0315_\[4\] _01703_ VPWR VGND sg13g2_nand3_1
Xhold1709 _01058_ VPWR VGND net3536 sg13g2_dlygate4sd3_1
X_09008__974 VPWR VGND net1394 sg13g2_tiehi
X_08547__109 VPWR VGND net109 sg13g2_tiehi
X_06710_ VPWR VGND _01506_ _02743_ _02744_ _01365_ _00662_ _02719_ sg13g2_a221oi_1
X_07690_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[25\]
+ net2727 net999 _01192_ VPWR VGND sg13g2_mux2_1
XFILLER_92_584 VPWR VGND sg13g2_fill_2
XFILLER_92_573 VPWR VGND sg13g2_fill_1
X_06641_ net2886 net1154 _02684_ VPWR VGND sg13g2_nor2_1
XFILLER_64_297 VPWR VGND sg13g2_fill_2
X_06572_ net3605 net1156 _02638_ VPWR VGND sg13g2_nor2_1
X_08311_ net367 VGND VPWR _00392_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[13\]
+ clknet_leaf_83_clk_regs sg13g2_dfrbpq_1
X_09291_ net1817 VGND VPWR _01346_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[17\]
+ clknet_leaf_177_clk_regs sg13g2_dfrbpq_1
X_05523_ _02212_ net3443 net1070 VPWR VGND sg13g2_nand2_1
X_08242_ net435 VGND VPWR net2219 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[9\]
+ clknet_leaf_57_clk_regs sg13g2_dfrbpq_1
X_05454_ _02136_ i_exotiny._1615_\[2\] _02137_ _02161_ VPWR VGND sg13g2_a21o_1
X_05385_ _02103_ _02104_ net3326 _02106_ VPWR VGND _02105_ sg13g2_nand4_1
X_08173_ net504 VGND VPWR net3350 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[4\]
+ clknet_leaf_110_clk_regs sg13g2_dfrbpq_1
X_09015__967 VPWR VGND net1387 sg13g2_tiehi
X_07124_ net1290 net1841 _00874_ VPWR VGND sg13g2_and2_1
X_07055_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[25\]
+ net2573 net1015 _00816_ VPWR VGND sg13g2_mux2_1
X_06006_ net2982 net877 _02493_ _02497_ VPWR VGND sg13g2_mux2_1
XFILLER_0_728 VPWR VGND sg13g2_decap_8
X_09061__921 VPWR VGND net1341 sg13g2_tiehi
XFILLER_101_133 VPWR VGND sg13g2_fill_2
X_07957_ net700 VGND VPWR net3401 i_exotiny.i_wb_spi.cnt_hbit_r\[2\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_1
X_06908_ VGND VPWR _01368_ _02908_ _00696_ _02906_ sg13g2_a21oi_1
X_07888_ net3150 net3066 net981 _01355_ VPWR VGND sg13g2_mux2_1
XFILLER_29_979 VPWR VGND sg13g2_fill_1
X_06839_ net2061 net1188 _02853_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_161_clk_regs clknet_5_7__leaf_clk_regs clknet_leaf_161_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_43_459 VPWR VGND sg13g2_fill_1
X_08509_ net171 VGND VPWR net2533 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[29\]
+ clknet_leaf_71_clk_regs sg13g2_dfrbpq_1
XFILLER_106_951 VPWR VGND sg13g2_decap_8
XFILLER_11_94 VPWR VGND sg13g2_fill_2
XFILLER_105_494 VPWR VGND sg13g2_decap_8
X_09177__805 VPWR VGND net805 sg13g2_tiehi
XFILLER_4_1002 VPWR VGND sg13g2_decap_8
XFILLER_74_540 VPWR VGND sg13g2_fill_1
XFILLER_46_220 VPWR VGND sg13g2_fill_1
XFILLER_61_201 VPWR VGND sg13g2_fill_1
XFILLER_34_415 VPWR VGND sg13g2_fill_2
XFILLER_46_264 VPWR VGND sg13g2_fill_2
XFILLER_46_275 VPWR VGND sg13g2_fill_2
XFILLER_50_908 VPWR VGND sg13g2_fill_1
XFILLER_36_91 VPWR VGND sg13g2_decap_8
XFILLER_43_960 VPWR VGND sg13g2_fill_2
XFILLER_15_684 VPWR VGND sg13g2_fill_1
Xinput11 uio_in[1] net11 VPWR VGND sg13g2_buf_2
XFILLER_30_698 VPWR VGND sg13g2_fill_2
X_08477__203 VPWR VGND net203 sg13g2_tiehi
X_08843__1143 VPWR VGND net1563 sg13g2_tiehi
X_05170_ _01898_ _01899_ net36 VPWR VGND sg13g2_nor2_1
Xhold828 _00997_ VPWR VGND net2655 sg13g2_dlygate4sd3_1
Xhold817 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[11\]
+ VPWR VGND net2644 sg13g2_dlygate4sd3_1
Xhold806 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[7\]
+ VPWR VGND net2633 sg13g2_dlygate4sd3_1
Xhold839 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[26\]
+ VPWR VGND net2666 sg13g2_dlygate4sd3_1
XFILLER_6_382 VPWR VGND sg13g2_fill_1
XFILLER_103_409 VPWR VGND sg13g2_decap_8
X_08197__480 VPWR VGND net480 sg13g2_tiehi
X_08860_ net1546 VGND VPWR net2957 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[27\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk VPWR VGND sg13g2_buf_8
X_09045__938 VPWR VGND net1358 sg13g2_tiehi
Xhold1506 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[13\]
+ VPWR VGND net3333 sg13g2_dlygate4sd3_1
X_07811_ net2680 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[29\]
+ net894 _01290_ VPWR VGND sg13g2_mux2_1
XFILLER_28_0 VPWR VGND sg13g2_decap_8
Xhold1517 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[7\]
+ VPWR VGND net3344 sg13g2_dlygate4sd3_1
Xhold1528 _00488_ VPWR VGND net3355 sg13g2_dlygate4sd3_1
Xhold1539 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[15\]
+ VPWR VGND net3366 sg13g2_dlygate4sd3_1
X_08791_ net1617 VGND VPWR _00849_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[22\]
+ clknet_leaf_169_clk_regs sg13g2_dfrbpq_1
X_07742_ _03207_ VPWR _03208_ VGND net2106 _03206_ sg13g2_o21ai_1
X_04954_ _01681_ _01682_ _01611_ _01686_ VPWR VGND _01685_ sg13g2_nand4_1
X_04885_ _01617_ net1258 net1260 VPWR VGND sg13g2_nand2_2
X_07673_ net2980 net3163 net1002 _01175_ VPWR VGND sg13g2_mux2_1
X_06624_ net1195 _02671_ _02672_ _00648_ VPWR VGND sg13g2_nor3_1
XFILLER_34_971 VPWR VGND sg13g2_fill_2
X_06555_ net1210 net3783 _02629_ _00622_ VPWR VGND sg13g2_a21o_1
XFILLER_33_470 VPWR VGND sg13g2_fill_2
X_06486_ net2876 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[13\]
+ net1025 _00567_ VPWR VGND sg13g2_mux2_1
X_09274_ net73 VGND VPWR net2070 i_exotiny._0021_\[0\] clknet_leaf_174_clk_regs sg13g2_dfrbpq_2
X_05506_ _02197_ VPWR i_exotiny._1611_\[15\] VGND net1074 _02199_ sg13g2_o21ai_1
X_05437_ net1232 _02133_ _02143_ _02146_ VPWR VGND sg13g2_nor3_1
X_08225_ net452 VGND VPWR net2710 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[24\]
+ clknet_leaf_170_clk_regs sg13g2_dfrbpq_1
X_08794__1194 VPWR VGND net1614 sg13g2_tiehi
X_05368_ _02082_ _02083_ _02079_ _02090_ VPWR VGND _02084_ sg13g2_nand4_1
X_08156_ net522 VGND VPWR net2258 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[20\]
+ clknet_leaf_132_clk_regs sg13g2_dfrbpq_1
XFILLER_4_319 VPWR VGND sg13g2_fill_2
X_07107_ net2216 _02945_ net914 _00858_ VPWR VGND sg13g2_mux2_1
XFILLER_106_7 VPWR VGND sg13g2_fill_1
X_08087_ net607 VGND VPWR _00168_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[24\]
+ clknet_leaf_86_clk_regs sg13g2_dfrbpq_1
X_05299_ VGND VPWR _02025_ i_exotiny._0018_\[0\] net1257 sg13g2_or2_1
XFILLER_106_258 VPWR VGND sg13g2_decap_8
X_07038_ net2548 net2410 net1013 _00799_ VPWR VGND sg13g2_mux2_1
XFILLER_102_420 VPWR VGND sg13g2_decap_8
XFILLER_103_965 VPWR VGND sg13g2_decap_8
XFILLER_88_687 VPWR VGND sg13g2_fill_2
X_08137__548 VPWR VGND net548 sg13g2_tiehi
XFILLER_102_497 VPWR VGND sg13g2_decap_8
XFILLER_75_337 VPWR VGND sg13g2_fill_2
X_08989_ net1413 VGND VPWR net2102 i_exotiny._1160_\[10\] clknet_leaf_164_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_84_860 VPWR VGND sg13g2_fill_1
XFILLER_56_573 VPWR VGND sg13g2_decap_8
X_08113__581 VPWR VGND net581 sg13g2_tiehi
XFILLER_43_278 VPWR VGND sg13g2_fill_2
XFILLER_7_168 VPWR VGND sg13g2_fill_2
XFILLER_4_820 VPWR VGND sg13g2_decap_8
XFILLER_99_919 VPWR VGND sg13g2_decap_8
XFILLER_98_418 VPWR VGND sg13g2_decap_8
X_08120__574 VPWR VGND net574 sg13g2_tiehi
XFILLER_4_897 VPWR VGND sg13g2_decap_8
XFILLER_105_291 VPWR VGND sg13g2_decap_8
Xfanout1120 _01582_ net1120 VPWR VGND sg13g2_buf_1
Xfanout1131 net1136 net1131 VPWR VGND sg13g2_buf_2
Xfanout1153 net1154 net1153 VPWR VGND sg13g2_buf_8
Xfanout1142 _02422_ net1142 VPWR VGND sg13g2_buf_8
Xfanout1164 _02414_ net1164 VPWR VGND sg13g2_buf_2
Xfanout1175 net1179 net1175 VPWR VGND sg13g2_buf_8
Xfanout1186 net1187 net1186 VPWR VGND sg13g2_buf_8
Xfanout1197 net1200 net1197 VPWR VGND sg13g2_buf_8
XFILLER_93_189 VPWR VGND sg13g2_fill_1
X_09005__977 VPWR VGND net1397 sg13g2_tiehi
X_04670_ net1242 net1245 net1247 _01431_ VPWR VGND sg13g2_nor3_2
XFILLER_47_595 VPWR VGND sg13g2_fill_2
XFILLER_90_896 VPWR VGND sg13g2_fill_1
XFILLER_50_727 VPWR VGND sg13g2_fill_1
X_06340_ net3044 net873 _02558_ _02563_ VPWR VGND sg13g2_mux2_1
X_09051__931 VPWR VGND net1351 sg13g2_tiehi
X_06271_ net2647 net2814 net943 _00414_ VPWR VGND sg13g2_mux2_1
XFILLER_30_473 VPWR VGND sg13g2_fill_2
X_08010_ net685 VGND VPWR _00091_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[11\]
+ clknet_leaf_61_clk_regs sg13g2_dfrbpq_1
X_05222_ _01947_ _01948_ _01946_ _01950_ VPWR VGND _01949_ sg13g2_nand4_1
Xhold603 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[31\]
+ VPWR VGND net2430 sg13g2_dlygate4sd3_1
Xhold636 _01137_ VPWR VGND net2463 sg13g2_dlygate4sd3_1
X_09229__750 VPWR VGND net750 sg13g2_tiehi
Xhold625 _01331_ VPWR VGND net2452 sg13g2_dlygate4sd3_1
Xhold614 _00183_ VPWR VGND net2441 sg13g2_dlygate4sd3_1
X_05153_ VGND VPWR i_exotiny._0043_\[2\] _01621_ _01883_ _01882_ sg13g2_a21oi_1
XFILLER_103_206 VPWR VGND sg13g2_decap_8
Xhold669 _01019_ VPWR VGND net2496 sg13g2_dlygate4sd3_1
Xhold647 _00496_ VPWR VGND net2474 sg13g2_dlygate4sd3_1
Xhold658 _00080_ VPWR VGND net2485 sg13g2_dlygate4sd3_1
X_05084_ _01677_ _01815_ net41 VPWR VGND sg13g2_nor2_1
XFILLER_98_930 VPWR VGND sg13g2_decap_8
X_08912_ net1490 VGND VPWR _00970_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[10\]
+ clknet_leaf_64_clk_regs sg13g2_dfrbpq_1
Xhold2015 i_exotiny.i_wdg_top.clk_div_inst.cnt\[15\] VPWR VGND net3842 sg13g2_dlygate4sd3_1
Xhold2004 i_exotiny._0077_\[4\] VPWR VGND net3831 sg13g2_dlygate4sd3_1
XFILLER_100_924 VPWR VGND sg13g2_decap_8
Xhold1325 _00546_ VPWR VGND net3152 sg13g2_dlygate4sd3_1
X_08843_ net1563 VGND VPWR net2788 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[10\]
+ clknet_leaf_185_clk_regs sg13g2_dfrbpq_1
Xhold1314 _01336_ VPWR VGND net3141 sg13g2_dlygate4sd3_1
Xhold1303 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[15\]
+ VPWR VGND net3130 sg13g2_dlygate4sd3_1
Xhold1347 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[31\]
+ VPWR VGND net3174 sg13g2_dlygate4sd3_1
X_05986_ net2154 net3234 net1050 _00188_ VPWR VGND sg13g2_mux2_1
Xhold1358 i_exotiny._0315_\[23\] VPWR VGND net3185 sg13g2_dlygate4sd3_1
X_08774_ net1634 VGND VPWR net3040 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[5\]
+ clknet_leaf_169_clk_regs sg13g2_dfrbpq_1
Xhold1336 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[12\]
+ VPWR VGND net3163 sg13g2_dlygate4sd3_1
X_08702__1286 VPWR VGND net1706 sg13g2_tiehi
X_07725_ net3453 net2642 net996 _01221_ VPWR VGND sg13g2_mux2_1
Xhold1369 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[19\]
+ VPWR VGND net3196 sg13g2_dlygate4sd3_1
X_04937_ _01669_ _01621_ i_exotiny._0043_\[3\] _01618_ i_exotiny._0031_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_07656_ net3085 _03189_ net899 _01163_ VPWR VGND sg13g2_mux2_1
X_04868_ _01597_ _01600_ _01477_ i_exotiny._1266_ VPWR VGND sg13g2_nand3_1
X_07587_ _03163_ net3843 net1913 _03159_ VPWR VGND sg13g2_and3_1
X_04799_ net3651 _01487_ net1282 _01547_ VPWR VGND sg13g2_nand3_1
X_06607_ i_exotiny._0314_\[15\] net1163 _02661_ VPWR VGND sg13g2_nor2_1
X_06538_ net2782 net2491 net930 _00613_ VPWR VGND sg13g2_mux2_1
X_09257_ net550 VGND VPWR _01312_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[15\]
+ clknet_leaf_129_clk_regs sg13g2_dfrbpq_1
X_08208_ net469 VGND VPWR _00289_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[7\]
+ clknet_leaf_151_clk_regs sg13g2_dfrbpq_1
XFILLER_21_484 VPWR VGND sg13g2_fill_2
X_06469_ i_exotiny._0039_\[3\] net873 _02608_ _02613_ VPWR VGND sg13g2_mux2_1
X_09188_ net793 VGND VPWR net3058 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[10\]
+ clknet_leaf_79_clk_regs sg13g2_dfrbpq_1
X_08924__1058 VPWR VGND net1478 sg13g2_tiehi
X_09167__815 VPWR VGND net815 sg13g2_tiehi
X_08139_ net546 VGND VPWR net2514 i_exotiny._0025_\[3\] clknet_leaf_118_clk_regs sg13g2_dfrbpq_2
XFILLER_104_4 VPWR VGND sg13g2_fill_1
XFILLER_1_845 VPWR VGND sg13g2_decap_8
XFILLER_103_762 VPWR VGND sg13g2_decap_8
XFILLER_89_974 VPWR VGND sg13g2_decap_8
XFILLER_48_304 VPWR VGND sg13g2_fill_1
XFILLER_102_294 VPWR VGND sg13g2_decap_8
X_08467__213 VPWR VGND net213 sg13g2_tiehi
Xhold1881 i_exotiny.i_wdg_top.o_wb_dat\[8\] VPWR VGND net3708 sg13g2_dlygate4sd3_1
Xhold1870 i_exotiny._1617_\[1\] VPWR VGND net3697 sg13g2_dlygate4sd3_1
XFILLER_72_830 VPWR VGND sg13g2_fill_1
XFILLER_57_893 VPWR VGND sg13g2_fill_2
X_09174__808 VPWR VGND net808 sg13g2_tiehi
XFILLER_1_1027 VPWR VGND sg13g2_fill_2
Xhold1892 i_exotiny._6090_\[2\] VPWR VGND net3719 sg13g2_dlygate4sd3_1
X_08187__490 VPWR VGND net490 sg13g2_tiehi
XFILLER_71_395 VPWR VGND sg13g2_fill_1
XFILLER_9_967 VPWR VGND sg13g2_decap_8
X_08474__206 VPWR VGND net206 sg13g2_tiehi
X_08194__483 VPWR VGND net483 sg13g2_tiehi
XFILLER_95_933 VPWR VGND sg13g2_decap_8
XFILLER_66_112 VPWR VGND sg13g2_fill_2
X_05840_ _02425_ _02426_ _01610_ _02429_ VPWR VGND _02427_ sg13g2_nand4_1
XFILLER_66_178 VPWR VGND sg13g2_fill_2
X_05771_ _02398_ i_exotiny._2034_\[4\] _00026_ VPWR VGND sg13g2_nand2_1
XFILLER_75_690 VPWR VGND sg13g2_decap_8
X_07510_ net3052 net3185 net904 _01093_ VPWR VGND sg13g2_mux2_1
X_08490_ net190 VGND VPWR _00564_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[10\]
+ clknet_leaf_94_clk_regs sg13g2_dfrbpq_1
X_04722_ VGND VPWR net1269 _01443_ _01480_ _01479_ sg13g2_a21oi_1
X_04653_ _01415_ net3777 VPWR VGND sg13g2_inv_2
X_07441_ net3307 net1215 _03083_ VPWR VGND sg13g2_and2_1
XFILLER_50_557 VPWR VGND sg13g2_fill_2
X_07372_ net3010 net1078 _03030_ VPWR VGND sg13g2_nor2_1
X_09111_ net871 VGND VPWR net3146 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[31\]
+ clknet_leaf_144_clk_regs sg13g2_dfrbpq_1
X_06323_ net2113 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[17\]
+ net1034 _00460_ VPWR VGND sg13g2_mux2_1
X_06254_ net2741 net2200 net1041 _00403_ VPWR VGND sg13g2_mux2_1
X_09042_ net1360 VGND VPWR _01100_ i_exotiny._0315_\[30\] clknet_leaf_2_clk_regs sg13g2_dfrbpq_2
X_06185_ net3161 _02537_ net952 _00344_ VPWR VGND sg13g2_mux2_1
Xhold400 _00335_ VPWR VGND net2227 sg13g2_dlygate4sd3_1
Xhold411 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[23\]
+ VPWR VGND net2238 sg13g2_dlygate4sd3_1
X_05205_ _01926_ _01931_ _01924_ _01933_ VPWR VGND _01932_ sg13g2_nand4_1
Xhold433 _01347_ VPWR VGND net2260 sg13g2_dlygate4sd3_1
Xhold444 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[30\]
+ VPWR VGND net2271 sg13g2_dlygate4sd3_1
Xhold422 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[29\]
+ VPWR VGND net2249 sg13g2_dlygate4sd3_1
X_05136_ VPWR VGND i_exotiny._0028_\[2\] _01865_ _01781_ i_exotiny._0030_\[2\] _01866_
+ _01766_ sg13g2_a221oi_1
XFILLER_104_537 VPWR VGND sg13g2_decap_8
Xhold466 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[9\]
+ VPWR VGND net2293 sg13g2_dlygate4sd3_1
Xhold477 _00253_ VPWR VGND net2304 sg13g2_dlygate4sd3_1
Xhold455 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[12\]
+ VPWR VGND net2282 sg13g2_dlygate4sd3_1
X_08103__591 VPWR VGND net591 sg13g2_tiehi
Xhold499 _00455_ VPWR VGND net2326 sg13g2_dlygate4sd3_1
Xfanout924 net928 net924 VPWR VGND sg13g2_buf_8
Xhold488 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[23\]
+ VPWR VGND net2315 sg13g2_dlygate4sd3_1
Xfanout913 net915 net913 VPWR VGND sg13g2_buf_8
Xfanout902 net903 net902 VPWR VGND sg13g2_buf_8
X_05067_ _01796_ _01797_ _01793_ _01799_ VPWR VGND _01798_ sg13g2_nand4_1
Xfanout968 net970 net968 VPWR VGND sg13g2_buf_8
Xfanout957 _02520_ net957 VPWR VGND sg13g2_buf_8
Xfanout946 net949 net946 VPWR VGND sg13g2_buf_8
Xhold1100 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[30\]
+ VPWR VGND net2927 sg13g2_dlygate4sd3_1
Xfanout935 net936 net935 VPWR VGND sg13g2_buf_8
X_08826_ net1582 VGND VPWR _00884_ i_exotiny.i_wb_spi.state_r\[25\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_86_966 VPWR VGND sg13g2_fill_1
Xfanout979 net980 net979 VPWR VGND sg13g2_buf_8
Xhold1122 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[22\]
+ VPWR VGND net2949 sg13g2_dlygate4sd3_1
Xhold1111 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[23\]
+ VPWR VGND net2938 sg13g2_dlygate4sd3_1
Xhold1133 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[15\]
+ VPWR VGND net2960 sg13g2_dlygate4sd3_1
XFILLER_46_808 VPWR VGND sg13g2_fill_2
XFILLER_100_765 VPWR VGND sg13g2_fill_2
Xhold1166 _01199_ VPWR VGND net2993 sg13g2_dlygate4sd3_1
Xhold1144 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[31\]
+ VPWR VGND net2971 sg13g2_dlygate4sd3_1
XFILLER_39_871 VPWR VGND sg13g2_fill_1
Xhold1155 i_exotiny._0013_\[2\] VPWR VGND net2982 sg13g2_dlygate4sd3_1
XFILLER_100_798 VPWR VGND sg13g2_fill_2
X_08757_ net1651 VGND VPWR net2831 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[20\]
+ clknet_leaf_80_clk_regs sg13g2_dfrbpq_1
X_05969_ i_exotiny._0020_\[3\] net874 _02486_ _02491_ VPWR VGND sg13g2_mux2_1
Xhold1199 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[6\]
+ VPWR VGND net3026 sg13g2_dlygate4sd3_1
Xhold1188 _00294_ VPWR VGND net3015 sg13g2_dlygate4sd3_1
Xhold1177 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[26\]
+ VPWR VGND net3004 sg13g2_dlygate4sd3_1
X_08688_ net1720 VGND VPWR net2281 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[15\]
+ clknet_leaf_105_clk_regs sg13g2_dfrbpq_1
XFILLER_54_863 VPWR VGND sg13g2_fill_1
X_07708_ net2545 net2959 net994 _01204_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_68_clk_regs clknet_5_24__leaf_clk_regs clknet_leaf_68_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_53_373 VPWR VGND sg13g2_fill_2
XFILLER_13_215 VPWR VGND sg13g2_fill_2
X_07639_ net2958 net2785 net899 _01147_ VPWR VGND sg13g2_mux2_1
XFILLER_53_395 VPWR VGND sg13g2_fill_1
X_08110__584 VPWR VGND net584 sg13g2_tiehi
XFILLER_16_1013 VPWR VGND sg13g2_fill_1
XFILLER_10_977 VPWR VGND sg13g2_decap_8
XFILLER_6_948 VPWR VGND sg13g2_decap_8
X_09273__75 VPWR VGND net75 sg13g2_tiehi
X_09180__801 VPWR VGND net801 sg13g2_tiehi
XFILLER_95_32 VPWR VGND sg13g2_fill_2
XFILLER_89_793 VPWR VGND sg13g2_fill_2
XFILLER_49_624 VPWR VGND sg13g2_fill_2
XFILLER_0_163 VPWR VGND sg13g2_fill_2
XFILLER_103_592 VPWR VGND sg13g2_fill_2
XFILLER_76_454 VPWR VGND sg13g2_fill_1
XFILLER_64_616 VPWR VGND sg13g2_fill_2
X_09041__941 VPWR VGND net1361 sg13g2_tiehi
XFILLER_63_148 VPWR VGND sg13g2_fill_2
X_09219__760 VPWR VGND net760 sg13g2_tiehi
XFILLER_44_373 VPWR VGND sg13g2_fill_1
XFILLER_99_535 VPWR VGND sg13g2_fill_1
X_09226__753 VPWR VGND net753 sg13g2_tiehi
X_07990_ net131 VGND VPWR i_exotiny._1611_\[23\] i_exotiny._0369_\[15\] clknet_leaf_14_clk_regs
+ sg13g2_dfrbpq_2
X_06941_ net2503 net2747 net924 _00720_ VPWR VGND sg13g2_mux2_1
X_08611_ net1785 VGND VPWR _00683_ i_exotiny._1617_\[3\] clknet_leaf_23_clk_regs sg13g2_dfrbpq_2
X_06872_ VGND VPWR i_exotiny._1618_\[0\] net1128 _02881_ _02880_ sg13g2_a21oi_1
XFILLER_10_0 VPWR VGND sg13g2_fill_1
XFILLER_39_156 VPWR VGND sg13g2_fill_2
XFILLER_94_284 VPWR VGND sg13g2_decap_8
X_05823_ net2501 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[15\]
+ net1054 _00095_ VPWR VGND sg13g2_mux2_1
X_05754_ _02387_ net3399 _02385_ VPWR VGND sg13g2_nand2b_1
X_08542_ net138 VGND VPWR net3240 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[30\]
+ clknet_leaf_183_clk_regs sg13g2_dfrbpq_1
X_09157__825 VPWR VGND net825 sg13g2_tiehi
XFILLER_91_980 VPWR VGND sg13g2_decap_8
X_08473_ net207 VGND VPWR net2250 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[25\]
+ clknet_leaf_163_clk_regs sg13g2_dfrbpq_1
X_04705_ _01423_ _01428_ _01463_ VPWR VGND sg13g2_and2_1
X_05685_ VGND VPWR i_exotiny._1616_\[1\] net1121 _02335_ _02334_ sg13g2_a21oi_1
X_07424_ i_exotiny._1160_\[18\] net1215 _03070_ VPWR VGND sg13g2_nor2_1
X_04636_ VPWR _01398_ i_exotiny._2034_\[0\] VGND sg13g2_inv_1
XFILLER_51_899 VPWR VGND sg13g2_fill_2
X_09233__746 VPWR VGND net746 sg13g2_tiehi
X_07355_ _03017_ _03015_ _03016_ net1207 net3010 VPWR VGND sg13g2_a22oi_1
X_07286_ net2789 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[15\]
+ net911 _01003_ VPWR VGND sg13g2_mux2_1
X_06306_ net3429 net3260 net1034 _00443_ VPWR VGND sg13g2_mux2_1
XFILLER_40_16 VPWR VGND sg13g2_fill_2
X_06237_ net2415 net2136 net1039 _00386_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_186_clk_regs clknet_5_0__leaf_clk_regs clknet_leaf_186_clk_regs VPWR
+ VGND sg13g2_buf_8
X_09025_ net1377 VGND VPWR net3546 i_exotiny._0315_\[13\] clknet_leaf_181_clk_regs
+ sg13g2_dfrbpq_1
X_08457__223 VPWR VGND net223 sg13g2_tiehi
XFILLER_3_907 VPWR VGND sg13g2_decap_8
XFILLER_105_846 VPWR VGND sg13g2_decap_8
X_06168_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[16\]
+ net2109 net953 _00330_ VPWR VGND sg13g2_mux2_1
Xhold241 _01001_ VPWR VGND net2068 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_115_clk_regs clknet_5_7__leaf_clk_regs clknet_leaf_115_clk_regs VPWR
+ VGND sg13g2_buf_8
Xhold252 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[7\]
+ VPWR VGND net2079 sg13g2_dlygate4sd3_1
X_09164__818 VPWR VGND net818 sg13g2_tiehi
Xhold230 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[11\]
+ VPWR VGND net2057 sg13g2_dlygate4sd3_1
XFILLER_104_334 VPWR VGND sg13g2_decap_8
Xhold296 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[22\]
+ VPWR VGND net2123 sg13g2_dlygate4sd3_1
X_06099_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[25\]
+ net2400 net955 _00275_ VPWR VGND sg13g2_mux2_1
Xhold285 _00785_ VPWR VGND net2112 sg13g2_dlygate4sd3_1
XFILLER_6_8 VPWR VGND sg13g2_decap_8
Xhold274 i_exotiny._1160_\[10\] VPWR VGND net2101 sg13g2_dlygate4sd3_1
X_05119_ _01849_ i_exotiny._0019_\[2\] _01773_ VPWR VGND sg13g2_nand2_1
Xhold263 _00768_ VPWR VGND net2090 sg13g2_dlygate4sd3_1
XFILLER_77_218 VPWR VGND sg13g2_fill_2
X_08856__1130 VPWR VGND net1550 sg13g2_tiehi
XFILLER_105_75 VPWR VGND sg13g2_decap_8
XFILLER_105_97 VPWR VGND sg13g2_fill_1
X_08809_ net1599 VGND VPWR _00867_ i_exotiny.i_wb_spi.state_r\[8\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_58_487 VPWR VGND sg13g2_fill_1
X_08464__216 VPWR VGND net216 sg13g2_tiehi
XFILLER_92_1026 VPWR VGND sg13g2_fill_2
X_08184__493 VPWR VGND net493 sg13g2_tiehi
XFILLER_6_734 VPWR VGND sg13g2_fill_1
XFILLER_5_266 VPWR VGND sg13g2_fill_2
X_08661__1316 VPWR VGND net1736 sg13g2_tiehi
X_08471__209 VPWR VGND net209 sg13g2_tiehi
X_08191__486 VPWR VGND net486 sg13g2_tiehi
XFILLER_65_914 VPWR VGND sg13g2_fill_1
Xinput9 ui_in[7] net9 VPWR VGND sg13g2_buf_1
XFILLER_36_104 VPWR VGND sg13g2_decap_4
XFILLER_91_221 VPWR VGND sg13g2_fill_1
X_05470_ i_exotiny._1611_\[1\] net1281 net3702 net11 VPWR VGND sg13g2_and3_1
X_07140_ net1286 net1854 _00890_ VPWR VGND sg13g2_and2_1
X_08556__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_69_1028 VPWR VGND sg13g2_fill_1
X_07071_ _02940_ net1142 net1163 _02941_ VPWR VGND sg13g2_a21o_1
XFILLER_105_109 VPWR VGND sg13g2_decap_8
X_06022_ VGND VPWR net3622 net1104 _00213_ _02505_ sg13g2_a21oi_1
XFILLER_99_332 VPWR VGND sg13g2_decap_8
X_08637__1340 VPWR VGND net1760 sg13g2_tiehi
XFILLER_59_229 VPWR VGND sg13g2_fill_1
X_08100__594 VPWR VGND net594 sg13g2_tiehi
X_07973_ net114 VGND VPWR i_exotiny._1611_\[1\] i_exotiny._0369_\[25\] clknet_leaf_10_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_101_359 VPWR VGND sg13g2_decap_8
XFILLER_56_903 VPWR VGND sg13g2_fill_2
X_06924_ net2635 net2688 net926 _00703_ VPWR VGND sg13g2_mux2_1
XFILLER_83_744 VPWR VGND sg13g2_fill_1
X_06855_ net3572 net1096 _02867_ VPWR VGND sg13g2_nor2_1
X_05806_ net1184 VPWR _02423_ VGND i_exotiny._1265_ net1162 sg13g2_o21ai_1
XFILLER_70_416 VPWR VGND sg13g2_fill_1
XFILLER_64_991 VPWR VGND sg13g2_fill_1
X_06786_ VGND VPWR net3630 net1133 _02809_ _02808_ sg13g2_a21oi_1
X_08525_ net155 VGND VPWR _00599_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[13\]
+ clknet_leaf_177_clk_regs sg13g2_dfrbpq_1
X_05737_ _02374_ net1118 _02372_ VPWR VGND sg13g2_nand2_1
XFILLER_23_321 VPWR VGND sg13g2_fill_1
X_05668_ net1123 i_exotiny._1924_\[17\] _02322_ VPWR VGND sg13g2_nor2b_1
X_08456_ net224 VGND VPWR net2610 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[8\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_1
XFILLER_51_663 VPWR VGND sg13g2_fill_2
X_07986__127 VPWR VGND net127 sg13g2_tiehi
X_08387_ net291 VGND VPWR net2731 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[25\]
+ clknet_leaf_139_clk_regs sg13g2_dfrbpq_1
X_04619_ VPWR _01381_ net3726 VGND sg13g2_inv_1
X_07407_ net1085 net2065 _03057_ _01046_ VPWR VGND sg13g2_a21o_1
X_05599_ VGND VPWR _01361_ net1105 _00024_ _02270_ sg13g2_a21oi_1
X_07338_ _02999_ _03001_ _03002_ VPWR VGND sg13g2_nor2_1
XFILLER_100_1008 VPWR VGND sg13g2_decap_8
X_07269_ i_exotiny._0040_\[2\] net880 _02972_ _02976_ VPWR VGND sg13g2_mux2_1
X_09031__951 VPWR VGND net1371 sg13g2_tiehi
X_09008_ net1394 VGND VPWR _01066_ i_exotiny._0079_\[1\] clknet_leaf_161_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_105_643 VPWR VGND sg13g2_decap_8
XFILLER_104_131 VPWR VGND sg13g2_decap_8
X_09209__770 VPWR VGND net770 sg13g2_tiehi
XFILLER_78_538 VPWR VGND sg13g2_decap_8
X_07947__94 VPWR VGND net94 sg13g2_tiehi
XFILLER_101_871 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_83_clk_regs clknet_5_27__leaf_clk_regs clknet_leaf_83_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_73_210 VPWR VGND sg13g2_fill_1
XFILLER_100_381 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_12_clk_regs clknet_5_3__leaf_clk_regs clknet_leaf_12_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_27_693 VPWR VGND sg13g2_fill_1
X_08679__1309 VPWR VGND net1729 sg13g2_tiehi
XFILLER_15_866 VPWR VGND sg13g2_fill_1
X_09216__763 VPWR VGND net763 sg13g2_tiehi
XFILLER_41_151 VPWR VGND sg13g2_fill_2
X_08715__1273 VPWR VGND net1693 sg13g2_tiehi
X_08610__1366 VPWR VGND net1786 sg13g2_tiehi
X_09147__835 VPWR VGND net835 sg13g2_tiehi
X_08937__1045 VPWR VGND net1465 sg13g2_tiehi
XFILLER_96_357 VPWR VGND sg13g2_decap_8
X_09223__756 VPWR VGND net756 sg13g2_tiehi
X_04970_ VPWR _01702_ _01701_ VGND sg13g2_inv_1
XFILLER_77_582 VPWR VGND sg13g2_fill_1
XFILLER_37_402 VPWR VGND sg13g2_fill_1
XFILLER_38_947 VPWR VGND sg13g2_fill_2
X_06640_ net1965 net1161 _02683_ VPWR VGND sg13g2_nor2_1
X_08447__233 VPWR VGND net233 sg13g2_tiehi
XFILLER_52_427 VPWR VGND sg13g2_fill_2
X_09154__828 VPWR VGND net828 sg13g2_tiehi
X_06571_ net3390 net1162 _02637_ VPWR VGND sg13g2_nor2_1
XFILLER_46_991 VPWR VGND sg13g2_fill_1
X_08310_ net368 VGND VPWR _00391_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[12\]
+ clknet_leaf_83_clk_regs sg13g2_dfrbpq_1
X_09290_ net1819 VGND VPWR net2328 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[16\]
+ clknet_leaf_175_clk_regs sg13g2_dfrbpq_1
X_05522_ _02209_ VPWR i_exotiny._1611_\[21\] VGND net1074 _02211_ sg13g2_o21ai_1
XFILLER_36_1005 VPWR VGND sg13g2_fill_2
X_08241_ net436 VGND VPWR net3192 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[8\]
+ clknet_leaf_56_clk_regs sg13g2_dfrbpq_1
X_05453_ _02154_ VPWR net28 VGND _02159_ _02160_ sg13g2_o21ai_1
X_09295__1389 VPWR VGND net1809 sg13g2_tiehi
X_09230__749 VPWR VGND net749 sg13g2_tiehi
X_05384_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set[0]
+ VPWR _02105_ VGND net1832 _02074_ sg13g2_o21ai_1
X_08172_ net505 VGND VPWR net2304 i_exotiny._0038_\[3\] clknet_leaf_69_clk_regs sg13g2_dfrbpq_2
X_07123_ net1290 net1835 _00873_ VPWR VGND sg13g2_and2_1
X_07054_ net2830 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[20\]
+ net1013 _00815_ VPWR VGND sg13g2_mux2_1
X_08454__226 VPWR VGND net226 sg13g2_tiehi
X_06005_ net2898 _02496_ net1048 _00205_ VPWR VGND sg13g2_mux2_1
XFILLER_82_1025 VPWR VGND sg13g2_decap_4
X_07956_ net703 VGND VPWR _00063_ i_exotiny.i_wb_spi.cnt_hbit_r\[1\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_101_178 VPWR VGND sg13g2_fill_2
X_06907_ net2570 net1263 net3241 _02908_ VPWR VGND sg13g2_nand3_1
XFILLER_68_593 VPWR VGND sg13g2_fill_1
XFILLER_46_15 VPWR VGND sg13g2_decap_8
XFILLER_83_530 VPWR VGND sg13g2_fill_1
X_07887_ net2810 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[29\]
+ net978 _01354_ VPWR VGND sg13g2_mux2_1
XFILLER_83_585 VPWR VGND sg13g2_fill_2
X_06838_ VGND VPWR net1097 _02851_ _00682_ _02852_ sg13g2_a21oi_1
X_06769_ _02794_ net1875 net1183 VPWR VGND sg13g2_nand2_1
X_08461__219 VPWR VGND net219 sg13g2_tiehi
XFILLER_36_490 VPWR VGND sg13g2_fill_2
X_08508_ net172 VGND VPWR _00582_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[28\]
+ clknet_leaf_109_clk_regs sg13g2_dfrbpq_1
XFILLER_51_460 VPWR VGND sg13g2_fill_1
XFILLER_12_847 VPWR VGND sg13g2_fill_1
X_08439_ net246 VGND VPWR net3760 i_exotiny._0369_\[0\] clknet_leaf_11_clk_regs sg13g2_dfrbpq_1
Xclkbuf_leaf_130_clk_regs clknet_5_20__leaf_clk_regs clknet_leaf_130_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08181__496 VPWR VGND net496 sg13g2_tiehi
XFILLER_106_930 VPWR VGND sg13g2_decap_8
XFILLER_105_473 VPWR VGND sg13g2_decap_8
XFILLER_78_379 VPWR VGND sg13g2_fill_2
XFILLER_98_1021 VPWR VGND sg13g2_decap_8
X_08546__110 VPWR VGND net110 sg13g2_tiehi
XFILLER_59_1005 VPWR VGND sg13g2_fill_2
XFILLER_28_991 VPWR VGND sg13g2_fill_1
X_07949__707 VPWR VGND net707 sg13g2_tiehi
XFILLER_99_7 VPWR VGND sg13g2_fill_1
Xinput12 uio_in[2] net12 VPWR VGND sg13g2_buf_2
XFILLER_11_880 VPWR VGND sg13g2_fill_2
Xhold807 _01170_ VPWR VGND net2634 sg13g2_dlygate4sd3_1
Xhold818 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[16\]
+ VPWR VGND net2645 sg13g2_dlygate4sd3_1
Xhold829 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[25\]
+ VPWR VGND net2656 sg13g2_dlygate4sd3_1
Xhold1507 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[14\]
+ VPWR VGND net3334 sg13g2_dlygate4sd3_1
X_08790_ net1618 VGND VPWR _00848_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[21\]
+ clknet_leaf_168_clk_regs sg13g2_dfrbpq_1
X_07810_ net3225 net3017 net893 _01289_ VPWR VGND sg13g2_mux2_1
Xhold1529 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[6\]
+ VPWR VGND net3356 sg13g2_dlygate4sd3_1
XFILLER_85_828 VPWR VGND sg13g2_fill_2
X_07741_ _03207_ net3805 _03206_ VPWR VGND sg13g2_nand2_1
Xhold1518 _00525_ VPWR VGND net3345 sg13g2_dlygate4sd3_1
X_04953_ _01685_ _01601_ _01684_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_733 VPWR VGND sg13g2_fill_2
XFILLER_53_725 VPWR VGND sg13g2_fill_1
XFILLER_53_703 VPWR VGND sg13g2_fill_2
X_09021__961 VPWR VGND net1381 sg13g2_tiehi
X_07672_ net2633 net2882 net1001 _01174_ VPWR VGND sg13g2_mux2_1
X_04884_ _01616_ i_exotiny._0077_\[3\] VPWR VGND i_exotiny._0077_\[2\] sg13g2_nand2b_2
XFILLER_93_894 VPWR VGND sg13g2_decap_8
X_06623_ net2038 net1152 _02672_ VPWR VGND sg13g2_nor2_1
X_08587__1390 VPWR VGND net1810 sg13g2_tiehi
X_06554_ net3641 net1213 _02629_ VPWR VGND sg13g2_and2_1
XFILLER_18_490 VPWR VGND sg13g2_fill_2
X_05505_ VGND VPWR i_exotiny._0314_\[7\] net1280 _02199_ _02198_ sg13g2_a21oi_1
X_06485_ net2448 net3022 net1026 _00566_ VPWR VGND sg13g2_mux2_1
X_09273_ net75 VGND VPWR _01328_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[31\]
+ clknet_leaf_131_clk_regs sg13g2_dfrbpq_1
X_05436_ _02142_ _02144_ _02145_ VPWR VGND sg13g2_nor2_1
X_08224_ net453 VGND VPWR net2334 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[23\]
+ clknet_leaf_150_clk_regs sg13g2_dfrbpq_1
X_05367_ _02081_ VPWR _02089_ VGND _00021_ i_exotiny._2034_\[7\] sg13g2_o21ai_1
X_08155_ net523 VGND VPWR net2019 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[19\]
+ clknet_leaf_119_clk_regs sg13g2_dfrbpq_1
XFILLER_10_1019 VPWR VGND sg13g2_decap_8
X_07106_ net3002 net872 _02940_ _02945_ VPWR VGND sg13g2_mux2_1
XFILLER_106_237 VPWR VGND sg13g2_decap_8
X_08086_ net608 VGND VPWR net2457 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[23\]
+ clknet_leaf_92_clk_regs sg13g2_dfrbpq_1
X_05298_ _02021_ _02022_ _02020_ _02024_ VPWR VGND _02023_ sg13g2_nand4_1
X_07037_ net3109 net3065 net1014 _00798_ VPWR VGND sg13g2_mux2_1
XFILLER_103_944 VPWR VGND sg13g2_decap_8
X_09206__773 VPWR VGND net773 sg13g2_tiehi
XFILLER_102_476 VPWR VGND sg13g2_decap_8
X_08988_ net1414 VGND VPWR net2066 i_exotiny._1160_\[9\] clknet_leaf_18_clk_regs sg13g2_dfrbpq_1
X_07939_ net709 VGND VPWR net1929 i_exotiny.i_wb_spi.spi_sdo_o clknet_leaf_29_clk_regs
+ sg13g2_dfrbpq_1
X_08629__774 VPWR VGND net774 sg13g2_tiehi
XFILLER_28_243 VPWR VGND sg13g2_fill_2
XFILLER_71_511 VPWR VGND sg13g2_fill_2
XFILLER_16_438 VPWR VGND sg13g2_fill_1
XFILLER_73_68 VPWR VGND sg13g2_fill_2
X_09137__845 VPWR VGND net845 sg13g2_tiehi
XFILLER_106_1014 VPWR VGND sg13g2_decap_8
XFILLER_89_1009 VPWR VGND sg13g2_decap_8
X_09213__766 VPWR VGND net766 sg13g2_tiehi
XFILLER_4_876 VPWR VGND sg13g2_decap_8
XFILLER_105_270 VPWR VGND sg13g2_decap_8
XFILLER_98_98 VPWR VGND sg13g2_fill_2
X_09144__838 VPWR VGND net838 sg13g2_tiehi
Xfanout1121 net1122 net1121 VPWR VGND sg13g2_buf_2
Xfanout1132 net1134 net1132 VPWR VGND sg13g2_buf_8
Xfanout1110 _01607_ net1110 VPWR VGND sg13g2_buf_8
Xfanout1143 _02390_ net1143 VPWR VGND sg13g2_buf_8
Xfanout1154 net1157 net1154 VPWR VGND sg13g2_buf_8
X_08566__72 VPWR VGND net72 sg13g2_tiehi
Xfanout1165 net1168 net1165 VPWR VGND sg13g2_buf_8
Xfanout1176 net1179 net1176 VPWR VGND sg13g2_buf_8
Xfanout1187 _01451_ net1187 VPWR VGND sg13g2_buf_8
X_09220__759 VPWR VGND net759 sg13g2_tiehi
Xfanout1198 net1199 net1198 VPWR VGND sg13g2_buf_8
XFILLER_47_563 VPWR VGND sg13g2_fill_1
XFILLER_62_555 VPWR VGND sg13g2_fill_1
X_08887__1095 VPWR VGND net1515 sg13g2_tiehi
X_06270_ net3026 i_exotiny._0016_\[2\] net939 _00413_ VPWR VGND sg13g2_mux2_1
X_05221_ _01949_ _01642_ i_exotiny._0015_\[1\] _01638_ i_exotiny._0029_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold604 _00143_ VPWR VGND net2431 sg13g2_dlygate4sd3_1
Xhold626 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[20\]
+ VPWR VGND net2453 sg13g2_dlygate4sd3_1
Xhold615 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[23\]
+ VPWR VGND net2442 sg13g2_dlygate4sd3_1
X_05152_ _01882_ _01873_ _01881_ VPWR VGND sg13g2_nand2_1
Xhold648 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[23\]
+ VPWR VGND net2475 sg13g2_dlygate4sd3_1
Xhold637 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[8\]
+ VPWR VGND net2464 sg13g2_dlygate4sd3_1
X_05083_ VPWR VGND _01814_ net1109 _01752_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[3\]
+ _01815_ net1107 sg13g2_a221oi_1
Xhold659 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[15\]
+ VPWR VGND net2486 sg13g2_dlygate4sd3_1
X_08911_ net1491 VGND VPWR _00969_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[9\]
+ clknet_leaf_112_clk_regs sg13g2_dfrbpq_1
X_08451__229 VPWR VGND net229 sg13g2_tiehi
XFILLER_40_0 VPWR VGND sg13g2_decap_4
XFILLER_100_903 VPWR VGND sg13g2_decap_8
XFILLER_97_452 VPWR VGND sg13g2_fill_1
Xhold2016 i_exotiny.i_wdg_top.clk_div_inst.cnt\[5\] VPWR VGND net3843 sg13g2_dlygate4sd3_1
Xhold2005 i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[1\] VPWR VGND net3832 sg13g2_dlygate4sd3_1
XFILLER_98_986 VPWR VGND sg13g2_decap_8
Xhold1304 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[14\]
+ VPWR VGND net3131 sg13g2_dlygate4sd3_1
Xhold1315 i_exotiny._1612_\[1\] VPWR VGND net3142 sg13g2_dlygate4sd3_1
XFILLER_69_176 VPWR VGND sg13g2_fill_1
X_08842_ net1564 VGND VPWR net2829 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[9\]
+ clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
Xhold1337 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[29\]
+ VPWR VGND net3164 sg13g2_dlygate4sd3_1
Xhold1359 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[13\]
+ VPWR VGND net3186 sg13g2_dlygate4sd3_1
X_08674__1314 VPWR VGND net1734 sg13g2_tiehi
Xhold1326 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[8\]
+ VPWR VGND net3153 sg13g2_dlygate4sd3_1
X_08773_ net1635 VGND VPWR net3001 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[4\]
+ clknet_leaf_168_clk_regs sg13g2_dfrbpq_1
XFILLER_38_530 VPWR VGND sg13g2_decap_8
Xhold1348 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[29\]
+ VPWR VGND net3175 sg13g2_dlygate4sd3_1
X_05985_ net2440 net2486 net1051 _00187_ VPWR VGND sg13g2_mux2_1
XFILLER_84_179 VPWR VGND sg13g2_fill_1
X_07724_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[25\]
+ net2748 net993 _01220_ VPWR VGND sg13g2_mux2_1
XFILLER_38_563 VPWR VGND sg13g2_fill_2
X_04936_ _01668_ _01655_ i_exotiny._0026_\[3\] _01642_ i_exotiny._0015_\[3\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_81_820 VPWR VGND sg13g2_fill_1
XFILLER_65_360 VPWR VGND sg13g2_fill_1
X_07655_ i_exotiny._0024_\[0\] net889 _03187_ _03189_ VPWR VGND sg13g2_mux2_1
X_06606_ net1199 _02659_ _02660_ _00642_ VPWR VGND sg13g2_nor3_1
X_04867_ VPWR VGND _01599_ _01454_ _01598_ net1269 _01600_ i_exotiny._1265_ sg13g2_a221oi_1
X_07586_ VGND VPWR i_exotiny.i_wdg_top.clk_div_inst.cnt\[5\] _03159_ _03162_ net1913
+ sg13g2_a21oi_1
X_04798_ net1283 VPWR _01546_ VGND i_exotiny._1623_ _01545_ sg13g2_o21ai_1
X_06537_ net2965 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[30\]
+ net929 _00612_ VPWR VGND sg13g2_mux2_1
X_06468_ _02612_ net3322 net937 _00552_ VPWR VGND sg13g2_mux2_1
X_09285__51 VPWR VGND net51 sg13g2_tiehi
X_09256_ net551 VGND VPWR _01311_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[14\]
+ clknet_leaf_126_clk_regs sg13g2_dfrbpq_1
X_05419_ _02127_ i_exotiny.i_wb_qspi_mem.cnt_r\[2\] _02128_ VPWR VGND sg13g2_xor2_1
X_08207_ net470 VGND VPWR _00288_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[6\]
+ clknet_leaf_152_clk_regs sg13g2_dfrbpq_1
X_08143__542 VPWR VGND net542 sg13g2_tiehi
X_09187_ net794 VGND VPWR net2901 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[9\]
+ clknet_leaf_80_clk_regs sg13g2_dfrbpq_1
X_08932__1050 VPWR VGND net1470 sg13g2_tiehi
X_06399_ _02574_ _02583_ _02584_ VPWR VGND sg13g2_nor2_1
X_08138_ net547 VGND VPWR _00219_ i_exotiny._0025_\[2\] clknet_leaf_118_clk_regs sg13g2_dfrbpq_2
X_08069_ net625 VGND VPWR _00150_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[6\]
+ clknet_leaf_86_clk_regs sg13g2_dfrbpq_1
XFILLER_1_824 VPWR VGND sg13g2_decap_8
XFILLER_103_741 VPWR VGND sg13g2_decap_8
XFILLER_89_953 VPWR VGND sg13g2_decap_8
XFILLER_102_273 VPWR VGND sg13g2_decap_8
Xhold1871 _02826_ VPWR VGND net3698 sg13g2_dlygate4sd3_1
Xhold1860 i_exotiny._1619_\[1\] VPWR VGND net3687 sg13g2_dlygate4sd3_1
XFILLER_1_1006 VPWR VGND sg13g2_decap_8
XFILLER_95_1024 VPWR VGND sg13g2_decap_4
Xhold1882 _02407_ VPWR VGND net3709 sg13g2_dlygate4sd3_1
XFILLER_17_736 VPWR VGND sg13g2_fill_1
Xhold1893 _00662_ VPWR VGND net3720 sg13g2_dlygate4sd3_1
XFILLER_72_875 VPWR VGND sg13g2_fill_1
X_08543__113 VPWR VGND net113 sg13g2_tiehi
XFILLER_17_769 VPWR VGND sg13g2_decap_4
XFILLER_9_946 VPWR VGND sg13g2_decap_8
XFILLER_13_997 VPWR VGND sg13g2_decap_8
X_08752__1236 VPWR VGND net1656 sg13g2_tiehi
X_09011__971 VPWR VGND net1391 sg13g2_tiehi
X_08550__106 VPWR VGND net106 sg13g2_tiehi
XFILLER_95_912 VPWR VGND sg13g2_decap_8
Xhold1 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[13\]
+ VPWR VGND net1828 sg13g2_dlygate4sd3_1
XFILLER_95_989 VPWR VGND sg13g2_decap_8
X_05770_ _02397_ VPWR _00069_ VGND net1143 _02396_ sg13g2_o21ai_1
X_04721_ net1174 _01471_ _01477_ _01479_ VPWR VGND sg13g2_nor3_1
X_08974__1008 VPWR VGND net1428 sg13g2_tiehi
X_04652_ VPWR _01414_ net1905 VGND sg13g2_inv_1
XFILLER_63_886 VPWR VGND sg13g2_fill_1
X_07440_ _03082_ VPWR _01054_ VGND net1083 _03081_ sg13g2_o21ai_1
X_07371_ _03029_ _03025_ _03028_ net1207 net2026 VPWR VGND sg13g2_a22oi_1
X_09110_ net1292 VGND VPWR net2297 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[30\]
+ clknet_leaf_143_clk_regs sg13g2_dfrbpq_1
X_06322_ net1976 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[16\]
+ net1035 _00459_ VPWR VGND sg13g2_mux2_1
X_09041_ net1361 VGND VPWR _01099_ i_exotiny._0315_\[29\] clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
X_06253_ net3159 net3357 net1038 _00402_ VPWR VGND sg13g2_mux2_1
X_06184_ net876 i_exotiny._0028_\[2\] _02533_ _02537_ VPWR VGND sg13g2_mux2_1
Xhold401 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[24\]
+ VPWR VGND net2228 sg13g2_dlygate4sd3_1
X_05204_ _01932_ _01783_ i_exotiny._0023_\[1\] _01767_ i_exotiny._0032_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold412 _00333_ VPWR VGND net2239 sg13g2_dlygate4sd3_1
X_08580__1402 VPWR VGND net1822 sg13g2_tiehi
Xhold434 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[22\]
+ VPWR VGND net2261 sg13g2_dlygate4sd3_1
Xhold445 _00243_ VPWR VGND net2272 sg13g2_dlygate4sd3_1
X_08728__1260 VPWR VGND net1680 sg13g2_tiehi
Xhold423 _00547_ VPWR VGND net2250 sg13g2_dlygate4sd3_1
X_05135_ _01863_ _01864_ _01862_ _01865_ VPWR VGND sg13g2_nand3_1
XFILLER_104_516 VPWR VGND sg13g2_decap_8
Xhold467 _00800_ VPWR VGND net2294 sg13g2_dlygate4sd3_1
Xhold456 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[14\]
+ VPWR VGND net2283 sg13g2_dlygate4sd3_1
Xhold478 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[29\]
+ VPWR VGND net2305 sg13g2_dlygate4sd3_1
Xfanout925 net928 net925 VPWR VGND sg13g2_buf_8
Xhold489 _00718_ VPWR VGND net2316 sg13g2_dlygate4sd3_1
X_09127__855 VPWR VGND net855 sg13g2_tiehi
Xfanout914 net915 net914 VPWR VGND sg13g2_buf_8
Xfanout903 net907 net903 VPWR VGND sg13g2_buf_8
X_05066_ _01798_ _01786_ i_exotiny._0017_\[3\] _01758_ i_exotiny._0040_\[3\] VPWR
+ VGND sg13g2_a22oi_1
Xfanout958 net959 net958 VPWR VGND sg13g2_buf_8
Xfanout947 net949 net947 VPWR VGND sg13g2_buf_8
Xfanout936 _02609_ net936 VPWR VGND sg13g2_buf_8
X_08825_ net1583 VGND VPWR _00883_ i_exotiny.i_wb_spi.state_r\[24\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_97_282 VPWR VGND sg13g2_decap_8
Xhold1112 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[19\]
+ VPWR VGND net2939 sg13g2_dlygate4sd3_1
Xfanout969 net971 net969 VPWR VGND sg13g2_buf_8
XFILLER_57_113 VPWR VGND sg13g2_fill_1
X_08623__1353 VPWR VGND net1773 sg13g2_tiehi
Xhold1123 _00461_ VPWR VGND net2950 sg13g2_dlygate4sd3_1
Xhold1101 _00725_ VPWR VGND net2928 sg13g2_dlygate4sd3_1
Xhold1156 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[5\]
+ VPWR VGND net2983 sg13g2_dlygate4sd3_1
Xhold1134 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[6\]
+ VPWR VGND net2961 sg13g2_dlygate4sd3_1
Xhold1145 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[11\]
+ VPWR VGND net2972 sg13g2_dlygate4sd3_1
Xhold1167 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[25\]
+ VPWR VGND net2994 sg13g2_dlygate4sd3_1
X_08756_ net1652 VGND VPWR net3426 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[19\]
+ clknet_leaf_87_clk_regs sg13g2_dfrbpq_1
X_05968_ net2477 _02490_ net967 _00174_ VPWR VGND sg13g2_mux2_1
Xhold1178 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[20\]
+ VPWR VGND net3005 sg13g2_dlygate4sd3_1
Xhold1189 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[19\]
+ VPWR VGND net3016 sg13g2_dlygate4sd3_1
XFILLER_26_522 VPWR VGND sg13g2_fill_1
X_05899_ net2482 net3092 net975 _00116_ VPWR VGND sg13g2_mux2_1
X_08687_ net1721 VGND VPWR net2330 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[14\]
+ clknet_leaf_104_clk_regs sg13g2_dfrbpq_1
X_04919_ net1256 _01620_ _01623_ _01651_ VPWR VGND sg13g2_nor3_2
X_07707_ net2990 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[4\]
+ net994 _01203_ VPWR VGND sg13g2_mux2_1
X_08830__1158 VPWR VGND net1578 sg13g2_tiehi
X_07638_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[11\]
+ net2706 net896 _01146_ VPWR VGND sg13g2_mux2_1
X_07902__48 VPWR VGND net48 sg13g2_tiehi
X_07569_ VGND VPWR net3699 net1231 _03152_ i_exotiny.i_wb_qspi_mem.cnt_r\[2\] sg13g2_a21oi_1
XFILLER_41_558 VPWR VGND sg13g2_decap_4
X_09134__848 VPWR VGND net848 sg13g2_tiehi
XFILLER_103_1028 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_37_clk_regs clknet_5_11__leaf_clk_regs clknet_leaf_37_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_10_956 VPWR VGND sg13g2_decap_8
XFILLER_6_927 VPWR VGND sg13g2_decap_8
X_09239_ net697 VGND VPWR net3376 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[29\]
+ clknet_leaf_130_clk_regs sg13g2_dfrbpq_1
X_09210__769 VPWR VGND net769 sg13g2_tiehi
Xhold990 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[10\]
+ VPWR VGND net2817 sg13g2_dlygate4sd3_1
XFILLER_62_1001 VPWR VGND sg13g2_fill_1
Xhold1690 i_exotiny._0314_\[11\] VPWR VGND net3517 sg13g2_dlygate4sd3_1
X_08480__200 VPWR VGND net200 sg13g2_tiehi
X_08806__1182 VPWR VGND net1602 sg13g2_tiehi
XFILLER_71_193 VPWR VGND sg13g2_fill_2
XFILLER_99_525 VPWR VGND sg13g2_fill_2
XFILLER_99_514 VPWR VGND sg13g2_decap_8
XFILLER_68_901 VPWR VGND sg13g2_fill_2
X_06940_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[20\]
+ net2192 net928 _00719_ VPWR VGND sg13g2_mux2_1
X_06871_ net1128 _02878_ _02879_ _02880_ VPWR VGND sg13g2_nor3_1
X_05822_ net2247 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[14\]
+ net1057 _00094_ VPWR VGND sg13g2_mux2_1
X_08610_ net1786 VGND VPWR net3564 i_exotiny._1617_\[2\] clknet_leaf_23_clk_regs sg13g2_dfrbpq_2
XFILLER_82_403 VPWR VGND sg13g2_fill_2
X_05753_ _01580_ _02386_ _00063_ VPWR VGND sg13g2_nor2_1
X_08541_ net139 VGND VPWR _00615_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[29\]
+ clknet_leaf_182_clk_regs sg13g2_dfrbpq_1
X_05684_ net1121 net1916 _02334_ VPWR VGND sg13g2_nor2b_1
X_08472_ net208 VGND VPWR net3152 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[24\]
+ clknet_leaf_64_clk_regs sg13g2_dfrbpq_1
X_04704_ _01462_ net1245 net1243 VPWR VGND sg13g2_nand2_1
X_04635_ VPWR _01397_ net1961 VGND sg13g2_inv_1
XFILLER_51_856 VPWR VGND sg13g2_fill_1
X_07423_ net1082 net2010 _03069_ _01050_ VPWR VGND sg13g2_a21o_1
XFILLER_50_355 VPWR VGND sg13g2_fill_2
X_07354_ net1207 _03013_ net1148 _03016_ VPWR VGND sg13g2_nor3_1
X_07285_ net2584 net2907 net909 _01002_ VPWR VGND sg13g2_mux2_1
X_06305_ VGND VPWR net1138 _02558_ _02559_ net1165 sg13g2_a21oi_1
X_06236_ net3087 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[6\]
+ net1038 _00385_ VPWR VGND sg13g2_mux2_1
X_09024_ net1378 VGND VPWR _01082_ i_exotiny._0315_\[12\] clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
Xhold220 _00048_ VPWR VGND net2047 sg13g2_dlygate4sd3_1
X_08140__545 VPWR VGND net545 sg13g2_tiehi
XFILLER_105_825 VPWR VGND sg13g2_decap_8
XFILLER_104_313 VPWR VGND sg13g2_decap_8
X_06167_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[15\]
+ net2263 net950 _00329_ VPWR VGND sg13g2_mux2_1
Xhold242 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[4\]
+ VPWR VGND net2069 sg13g2_dlygate4sd3_1
Xhold253 _00894_ VPWR VGND net2080 sg13g2_dlygate4sd3_1
Xhold231 _00529_ VPWR VGND net2058 sg13g2_dlygate4sd3_1
Xhold264 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[31\]
+ VPWR VGND net2091 sg13g2_dlygate4sd3_1
X_06098_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[24\]
+ net2276 net957 _00274_ VPWR VGND sg13g2_mux2_1
Xhold286 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[21\]
+ VPWR VGND net2113 sg13g2_dlygate4sd3_1
Xhold275 _01047_ VPWR VGND net2102 sg13g2_dlygate4sd3_1
X_05118_ _01848_ _01783_ i_exotiny._0023_\[2\] _01776_ i_exotiny._0021_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold297 _00130_ VPWR VGND net2124 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_155_clk_regs clknet_5_19__leaf_clk_regs clknet_leaf_155_clk_regs VPWR
+ VGND sg13g2_buf_8
X_05049_ net1238 net1240 net1220 _01781_ VGND VPWR _01759_ sg13g2_nor4_2
XFILLER_58_422 VPWR VGND sg13g2_fill_1
X_08808_ net1600 VGND VPWR _00866_ i_exotiny.i_wb_spi.state_r\[7\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_45_116 VPWR VGND sg13g2_fill_1
XFILLER_46_628 VPWR VGND sg13g2_fill_1
X_08739_ net1669 VGND VPWR _00797_ i_exotiny._0017_\[2\] clknet_leaf_84_clk_regs sg13g2_dfrbpq_2
XFILLER_73_469 VPWR VGND sg13g2_decap_4
XFILLER_92_1005 VPWR VGND sg13g2_decap_8
X_09001__981 VPWR VGND net1401 sg13g2_tiehi
XFILLER_30_61 VPWR VGND sg13g2_fill_2
XFILLER_30_94 VPWR VGND sg13g2_fill_2
XFILLER_2_985 VPWR VGND sg13g2_decap_8
XFILLER_17_374 VPWR VGND sg13g2_fill_2
XFILLER_33_867 VPWR VGND sg13g2_fill_1
X_09117__865 VPWR VGND net865 sg13g2_tiehi
X_07070_ _02420_ _02517_ _02940_ VPWR VGND sg13g2_nor2_2
X_06021_ net1888 net1104 _02505_ VPWR VGND sg13g2_nor2_1
XFILLER_99_311 VPWR VGND sg13g2_decap_8
XFILLER_99_388 VPWR VGND sg13g2_decap_8
XFILLER_102_839 VPWR VGND sg13g2_decap_8
XFILLER_101_338 VPWR VGND sg13g2_decap_8
X_07972_ net1178 VGND VPWR net1874 i_exotiny.i_wdg_top.o_wb_dat\[13\] clknet_leaf_58_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_56_915 VPWR VGND sg13g2_fill_2
X_06923_ net2720 net2721 net927 _00702_ VPWR VGND sg13g2_mux2_1
X_09124__858 VPWR VGND net858 sg13g2_tiehi
X_06854_ VGND VPWR i_exotiny._1619_\[1\] net1131 _02866_ _02865_ sg13g2_a21oi_1
XFILLER_28_628 VPWR VGND sg13g2_fill_1
XFILLER_71_907 VPWR VGND sg13g2_fill_1
X_06785_ net1132 _02806_ _02807_ _02808_ VPWR VGND sg13g2_nor3_1
X_05805_ VGND VPWR _01443_ net1157 _02422_ _01473_ sg13g2_a21oi_1
X_05736_ net1118 _02372_ _02373_ VPWR VGND sg13g2_and2_1
X_08524_ net156 VGND VPWR net2875 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[12\]
+ clknet_leaf_176_clk_regs sg13g2_dfrbpq_1
X_05667_ net1901 net1062 _02321_ VPWR VGND sg13g2_nor2_1
XFILLER_51_642 VPWR VGND sg13g2_decap_8
X_09170__812 VPWR VGND net812 sg13g2_tiehi
XFILLER_24_889 VPWR VGND sg13g2_fill_1
X_08455_ net225 VGND VPWR net2058 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[7\]
+ clknet_leaf_157_clk_regs sg13g2_dfrbpq_1
X_05598_ net3326 net1105 _02270_ VPWR VGND sg13g2_nor2_1
XFILLER_50_163 VPWR VGND sg13g2_fill_1
X_08386_ net292 VGND VPWR _00467_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[24\]
+ clknet_leaf_139_clk_regs sg13g2_dfrbpq_1
X_04618_ VPWR _01380_ net1270 VGND sg13g2_inv_1
X_07406_ net1085 _03055_ _03056_ _03057_ VPWR VGND sg13g2_nor3_1
X_07337_ VPWR _03001_ _03000_ VGND sg13g2_inv_1
X_07268_ _02975_ net2398 net1005 _00989_ VPWR VGND sg13g2_mux2_1
X_07199_ VGND VPWR _01409_ net1092 _00934_ _02961_ sg13g2_a21oi_1
X_06219_ net3208 net2717 net947 _00374_ VPWR VGND sg13g2_mux2_1
X_09007_ net1395 VGND VPWR _01065_ i_exotiny._0079_\[0\] clknet_leaf_160_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_105_622 VPWR VGND sg13g2_decap_8
X_08470__210 VPWR VGND net210 sg13g2_tiehi
XFILLER_2_226 VPWR VGND sg13g2_fill_1
XFILLER_105_699 VPWR VGND sg13g2_decap_8
XFILLER_104_187 VPWR VGND sg13g2_decap_8
XFILLER_101_850 VPWR VGND sg13g2_decap_8
XFILLER_100_360 VPWR VGND sg13g2_decap_8
XFILLER_19_639 VPWR VGND sg13g2_fill_2
XFILLER_33_119 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_52_clk_regs clknet_5_15__leaf_clk_regs clknet_leaf_52_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08687__1301 VPWR VGND net1721 sg13g2_tiehi
XFILLER_6_554 VPWR VGND sg13g2_fill_1
XFILLER_41_93 VPWR VGND sg13g2_fill_2
XFILLER_96_336 VPWR VGND sg13g2_decap_8
XFILLER_2_782 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_64_211 VPWR VGND sg13g2_fill_2
XFILLER_37_425 VPWR VGND sg13g2_fill_2
XFILLER_92_586 VPWR VGND sg13g2_fill_1
X_06570_ net1200 _02635_ _02636_ _00630_ VPWR VGND sg13g2_nor3_1
X_05521_ VGND VPWR i_exotiny._0314_\[13\] net1275 _02211_ _02210_ sg13g2_a21oi_1
XFILLER_33_653 VPWR VGND sg13g2_fill_1
X_08240_ net437 VGND VPWR _00321_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[7\]
+ clknet_leaf_60_clk_regs sg13g2_dfrbpq_1
X_05452_ net1264 VPWR _02160_ VGND i_exotiny._1619_\[1\] _02138_ sg13g2_o21ai_1
X_08171_ net506 VGND VPWR net2256 i_exotiny._0038_\[2\] clknet_leaf_70_clk_regs sg13g2_dfrbpq_2
X_08847__1139 VPWR VGND net1559 sg13g2_tiehi
XFILLER_21_848 VPWR VGND sg13g2_fill_2
X_07122_ net1289 net1837 _00872_ VPWR VGND sg13g2_and2_1
X_05383_ _02104_ _02073_ _02093_ VPWR VGND sg13g2_nand2_1
XFILLER_106_419 VPWR VGND sg13g2_decap_8
X_07053_ net3425 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[19\]
+ net1015 _00814_ VPWR VGND sg13g2_mux2_1
X_06004_ net2946 net882 _02493_ _02496_ VPWR VGND sg13g2_mux2_1
XFILLER_82_1004 VPWR VGND sg13g2_decap_8
XFILLER_87_325 VPWR VGND sg13g2_fill_2
XFILLER_102_658 VPWR VGND sg13g2_fill_2
X_07955_ net705 VGND VPWR _00062_ i_exotiny._1956_ clknet_leaf_32_clk_regs sg13g2_dfrbpq_2
X_08765__1223 VPWR VGND net1643 sg13g2_tiehi
X_06906_ _02907_ net2570 net1263 VPWR VGND sg13g2_nand2_1
XFILLER_56_701 VPWR VGND sg13g2_fill_2
X_07886_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[24\]
+ net2253 net979 _01353_ VPWR VGND sg13g2_mux2_1
X_06837_ net3563 net1097 _02852_ VPWR VGND sg13g2_nor2_1
X_06768_ VGND VPWR net1100 _02792_ _00671_ _02793_ sg13g2_a21oi_1
XFILLER_55_299 VPWR VGND sg13g2_fill_2
X_08507_ net173 VGND VPWR net2364 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[27\]
+ clknet_leaf_109_clk_regs sg13g2_dfrbpq_1
X_05719_ net1959 net1058 _02360_ VPWR VGND sg13g2_nor2_1
X_06699_ _02732_ _02734_ net1219 _02735_ VPWR VGND sg13g2_nand3_1
X_08438_ net247 VGND VPWR net3779 i_exotiny._0369_\[12\] clknet_leaf_16_clk_regs sg13g2_dfrbpq_2
X_08369_ net309 VGND VPWR _00450_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[7\]
+ clknet_leaf_133_clk_regs sg13g2_dfrbpq_1
XFILLER_20_870 VPWR VGND sg13g2_fill_2
XFILLER_20_892 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_170_clk_regs clknet_5_5__leaf_clk_regs clknet_leaf_170_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_106_986 VPWR VGND sg13g2_decap_8
XFILLER_105_452 VPWR VGND sg13g2_decap_8
XFILLER_11_96 VPWR VGND sg13g2_fill_1
XFILLER_98_1000 VPWR VGND sg13g2_decap_8
XFILLER_93_317 VPWR VGND sg13g2_decap_4
X_09107__875 VPWR VGND net1295 sg13g2_tiehi
XFILLER_93_339 VPWR VGND sg13g2_fill_2
XFILLER_47_789 VPWR VGND sg13g2_fill_1
XFILLER_46_277 VPWR VGND sg13g2_fill_1
XFILLER_43_940 VPWR VGND sg13g2_fill_1
Xinput13 uio_in[3] net13 VPWR VGND sg13g2_buf_2
X_09114__868 VPWR VGND net868 sg13g2_tiehi
XFILLER_7_852 VPWR VGND sg13g2_fill_2
Xhold808 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[4\]
+ VPWR VGND net2635 sg13g2_dlygate4sd3_1
Xhold819 _00779_ VPWR VGND net2646 sg13g2_dlygate4sd3_1
XFILLER_97_656 VPWR VGND sg13g2_fill_1
X_09160__822 VPWR VGND net822 sg13g2_tiehi
Xhold1508 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[8\]
+ VPWR VGND net3335 sg13g2_dlygate4sd3_1
X_07740_ net1119 _02946_ _03206_ VPWR VGND sg13g2_nor2_1
Xhold1519 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[31\]
+ VPWR VGND net3346 sg13g2_dlygate4sd3_1
X_04952_ _01684_ _01462_ _01463_ _01429_ _01427_ VPWR VGND sg13g2_a22oi_1
X_04883_ _01613_ _01614_ _01615_ VPWR VGND sg13g2_nor2_2
X_07671_ net2899 net3062 net1001 _01173_ VPWR VGND sg13g2_mux2_1
XFILLER_37_255 VPWR VGND sg13g2_fill_2
X_06622_ i_exotiny._0314_\[20\] net1159 _02671_ VPWR VGND sg13g2_nor2_1
X_06553_ net1210 net3794 _02628_ _00621_ VPWR VGND sg13g2_a21o_1
X_08460__220 VPWR VGND net220 sg13g2_tiehi
X_05504_ net1280 i_exotiny._0315_\[7\] _02198_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_472 VPWR VGND sg13g2_fill_1
XFILLER_34_973 VPWR VGND sg13g2_fill_1
XFILLER_34_984 VPWR VGND sg13g2_fill_1
X_06484_ net3195 net2578 net1023 _00565_ VPWR VGND sg13g2_mux2_1
X_09272_ net77 VGND VPWR _01327_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[30\]
+ clknet_leaf_123_clk_regs sg13g2_dfrbpq_1
X_05435_ _02144_ net1232 _02134_ VPWR VGND sg13g2_nand2_1
X_08223_ net454 VGND VPWR _00304_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[22\]
+ clknet_leaf_170_clk_regs sg13g2_dfrbpq_1
X_05366_ _02085_ _02086_ _02077_ _02088_ VPWR VGND _02087_ sg13g2_nand4_1
X_08154_ net524 VGND VPWR _00235_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[18\]
+ clknet_leaf_132_clk_regs sg13g2_dfrbpq_1
X_08085_ net609 VGND VPWR _00166_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[22\]
+ clknet_leaf_87_clk_regs sg13g2_dfrbpq_1
X_07105_ net3507 _02944_ net916 _00857_ VPWR VGND sg13g2_mux2_1
XFILLER_106_216 VPWR VGND sg13g2_decap_8
X_07036_ net3356 net2866 net1017 _00797_ VPWR VGND sg13g2_mux2_1
X_05297_ _02023_ _01632_ i_exotiny._0022_\[0\] _01622_ i_exotiny._0023_\[0\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_103_923 VPWR VGND sg13g2_decap_8
XFILLER_102_455 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_clk_regs clknet_0_clk_regs clknet_4_3_0_clk_regs VPWR VGND sg13g2_buf_8
X_08987_ net1415 VGND VPWR net2023 i_exotiny._1160_\[8\] clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
X_07938_ net710 VGND VPWR net1960 i_exotiny._1924_\[31\] clknet_leaf_30_clk_regs sg13g2_dfrbpq_1
X_07869_ net3140 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[11\]
+ net981 _01336_ VPWR VGND sg13g2_mux2_1
XFILLER_28_299 VPWR VGND sg13g2_fill_2
XFILLER_19_1001 VPWR VGND sg13g2_fill_1
XFILLER_4_855 VPWR VGND sg13g2_decap_8
XFILLER_106_783 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
Xfanout1111 _01577_ net1111 VPWR VGND sg13g2_buf_8
Xfanout1100 net1101 net1100 VPWR VGND sg13g2_buf_8
Xfanout1122 net1123 net1122 VPWR VGND sg13g2_buf_8
Xfanout1144 net1145 net1144 VPWR VGND sg13g2_buf_8
Xfanout1133 net1134 net1133 VPWR VGND sg13g2_buf_1
Xfanout1155 net1156 net1155 VPWR VGND sg13g2_buf_8
Xfanout1177 net1178 net1177 VPWR VGND sg13g2_buf_8
XFILLER_78_199 VPWR VGND sg13g2_fill_2
Xfanout1188 net1189 net1188 VPWR VGND sg13g2_buf_2
Xfanout1166 net1168 net1166 VPWR VGND sg13g2_buf_8
Xfanout1199 net1200 net1199 VPWR VGND sg13g2_buf_8
XFILLER_47_520 VPWR VGND sg13g2_fill_1
XFILLER_93_158 VPWR VGND sg13g2_fill_2
XFILLER_75_873 VPWR VGND sg13g2_fill_2
XFILLER_15_461 VPWR VGND sg13g2_fill_1
XFILLER_42_280 VPWR VGND sg13g2_fill_1
X_05220_ _01948_ _01653_ i_exotiny._0038_\[1\] _01618_ i_exotiny._0031_\[1\] VPWR
+ VGND sg13g2_a22oi_1
X_05151_ _01881_ _01628_ i_exotiny._0037_\[2\] _01624_ i_exotiny._0040_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold605 i_exotiny.i_wb_spi.dat_rx_r\[15\] VPWR VGND net2432 sg13g2_dlygate4sd3_1
Xhold627 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[23\]
+ VPWR VGND net2454 sg13g2_dlygate4sd3_1
Xhold616 _00914_ VPWR VGND net2443 sg13g2_dlygate4sd3_1
Xhold649 _00366_ VPWR VGND net2476 sg13g2_dlygate4sd3_1
Xhold638 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[5\]
+ VPWR VGND net2465 sg13g2_dlygate4sd3_1
X_05082_ VGND VPWR _01750_ _01813_ _01814_ net1108 sg13g2_a21oi_1
X_08910_ net1492 VGND VPWR net2879 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[8\]
+ clknet_leaf_65_clk_regs sg13g2_dfrbpq_1
Xhold2017 i_exotiny.i_wdg_top.clk_div_inst.cnt\[2\] VPWR VGND net3844 sg13g2_dlygate4sd3_1
XFILLER_98_965 VPWR VGND sg13g2_decap_8
Xhold2006 i_exotiny._1737_ VPWR VGND net3833 sg13g2_dlygate4sd3_1
X_08841_ net1565 VGND VPWR net2653 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[8\]
+ clknet_leaf_184_clk_regs sg13g2_dfrbpq_1
XFILLER_33_0 VPWR VGND sg13g2_decap_4
Xhold1316 _00208_ VPWR VGND net3143 sg13g2_dlygate4sd3_1
Xhold1305 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[13\]
+ VPWR VGND net3132 sg13g2_dlygate4sd3_1
XFILLER_100_959 VPWR VGND sg13g2_decap_8
Xhold1338 _00408_ VPWR VGND net3165 sg13g2_dlygate4sd3_1
X_05984_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[10\]
+ net2377 net1048 _00186_ VPWR VGND sg13g2_mux2_1
Xhold1327 _00594_ VPWR VGND net3154 sg13g2_dlygate4sd3_1
Xhold1349 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[11\]
+ VPWR VGND net3176 sg13g2_dlygate4sd3_1
X_08772_ net1636 VGND VPWR net2360 i_exotiny._0015_\[3\] clknet_leaf_163_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_72_309 VPWR VGND sg13g2_fill_2
X_07723_ net2048 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[20\]
+ net993 _01219_ VPWR VGND sg13g2_mux2_1
XFILLER_27_29 VPWR VGND sg13g2_fill_2
X_04935_ _01667_ _01641_ i_exotiny._0035_\[3\] _01615_ i_exotiny._0021_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_07654_ net2349 net3145 net896 _01162_ VPWR VGND sg13g2_mux2_1
XFILLER_26_748 VPWR VGND sg13g2_fill_2
X_06605_ net3402 net1156 _02660_ VPWR VGND sg13g2_nor2_1
X_04866_ net1270 net1267 _01599_ VPWR VGND sg13g2_nor2_1
X_07585_ net1204 _03161_ _01120_ VPWR VGND sg13g2_nor2_1
X_04797_ _01519_ i_exotiny._1757_ _01545_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_109_clk_regs clknet_5_28__leaf_clk_regs clknet_leaf_109_clk_regs VPWR
+ VGND sg13g2_buf_8
X_06536_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[25\]
+ net2150 net931 _00611_ VPWR VGND sg13g2_mux2_1
X_06467_ net3291 net877 _02608_ _02612_ VPWR VGND sg13g2_mux2_1
X_09255_ net552 VGND VPWR _01310_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[13\]
+ clknet_leaf_128_clk_regs sg13g2_dfrbpq_1
X_05418_ _01536_ _02126_ net1146 _02127_ VPWR VGND sg13g2_nand3_1
X_08206_ net471 VGND VPWR _00287_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[5\]
+ clknet_leaf_152_clk_regs sg13g2_dfrbpq_1
X_09186_ net795 VGND VPWR net2405 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[8\]
+ clknet_leaf_78_clk_regs sg13g2_dfrbpq_1
XFILLER_88_1021 VPWR VGND sg13g2_decap_8
X_06398_ net3665 net3509 net1272 _02583_ VPWR VGND sg13g2_mux2_1
X_05349_ i_exotiny.gpo\[0\] _02071_ gpo VPWR VGND sg13g2_and2_1
X_08137_ net548 VGND VPWR net3486 i_exotiny._0025_\[1\] clknet_leaf_132_clk_regs sg13g2_dfrbpq_2
X_08068_ net626 VGND VPWR net2419 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[5\]
+ clknet_leaf_93_clk_regs sg13g2_dfrbpq_1
XFILLER_103_720 VPWR VGND sg13g2_decap_8
XFILLER_1_803 VPWR VGND sg13g2_decap_8
X_07019_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[23\]
+ net3183 net918 _00786_ VPWR VGND sg13g2_mux2_1
XFILLER_102_252 VPWR VGND sg13g2_decap_8
XFILLER_103_797 VPWR VGND sg13g2_decap_8
Xhold1872 i_exotiny.i_wb_qspi_mem.cnt_r\[1\] VPWR VGND net3699 sg13g2_dlygate4sd3_1
Xhold1861 i_exotiny._0327_\[1\] VPWR VGND net3688 sg13g2_dlygate4sd3_1
X_09104__878 VPWR VGND net1298 sg13g2_tiehi
Xhold1850 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[1\] VPWR
+ VGND net3677 sg13g2_dlygate4sd3_1
XFILLER_95_1003 VPWR VGND sg13g2_decap_8
Xhold1883 _00074_ VPWR VGND net3710 sg13g2_dlygate4sd3_1
Xhold1894 i_exotiny.i_wb_regs.spi_size_o\[1\] VPWR VGND net3721 sg13g2_dlygate4sd3_1
X_08842__1144 VPWR VGND net1564 sg13g2_tiehi
XFILLER_17_40 VPWR VGND sg13g2_fill_2
X_09297__1349 VPWR VGND net1769 sg13g2_tiehi
XFILLER_9_925 VPWR VGND sg13g2_decap_8
X_09150__832 VPWR VGND net832 sg13g2_tiehi
XFILLER_13_976 VPWR VGND sg13g2_decap_8
XFILLER_24_291 VPWR VGND sg13g2_fill_2
XFILLER_106_580 VPWR VGND sg13g2_decap_8
X_08450__230 VPWR VGND net230 sg13g2_tiehi
XFILLER_95_968 VPWR VGND sg13g2_decap_8
Xhold2 _00804_ VPWR VGND net1829 sg13g2_dlygate4sd3_1
X_08793__1195 VPWR VGND net1615 sg13g2_tiehi
X_04720_ _01478_ _01477_ VPWR VGND sg13g2_inv_2
XFILLER_62_342 VPWR VGND sg13g2_fill_2
X_08982__1000 VPWR VGND net1420 sg13g2_tiehi
X_04651_ VPWR _01413_ net1897 VGND sg13g2_inv_1
XFILLER_35_567 VPWR VGND sg13g2_fill_1
X_07370_ net1872 net1217 _03028_ VPWR VGND sg13g2_and2_1
X_06321_ net3266 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[15\]
+ net1036 _00458_ VPWR VGND sg13g2_mux2_1
X_06252_ net2915 net2180 net1038 _00401_ VPWR VGND sg13g2_mux2_1
X_09040_ net1362 VGND VPWR net2100 i_exotiny._0315_\[28\] clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
X_05203_ _01931_ _01774_ i_exotiny._0018_\[1\] _01771_ i_exotiny._0016_\[1\] VPWR
+ VGND sg13g2_a22oi_1
X_06183_ net3023 _02536_ net951 _00343_ VPWR VGND sg13g2_mux2_1
Xhold402 _00574_ VPWR VGND net2229 sg13g2_dlygate4sd3_1
Xhold424 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[15\]
+ VPWR VGND net2251 sg13g2_dlygate4sd3_1
Xhold435 _00300_ VPWR VGND net2262 sg13g2_dlygate4sd3_1
Xhold413 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[12\]
+ VPWR VGND net2240 sg13g2_dlygate4sd3_1
X_05134_ _01864_ _01791_ i_exotiny._0026_\[2\] _01785_ i_exotiny._0043_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold457 _00485_ VPWR VGND net2284 sg13g2_dlygate4sd3_1
Xhold468 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[21\]
+ VPWR VGND net2295 sg13g2_dlygate4sd3_1
X_05065_ _01797_ _01783_ i_exotiny._0023_\[3\] _01782_ i_exotiny._0037_\[3\] VPWR
+ VGND sg13g2_a22oi_1
Xhold446 i_exotiny._0022_\[2\] VPWR VGND net2273 sg13g2_dlygate4sd3_1
Xhold479 _00372_ VPWR VGND net2306 sg13g2_dlygate4sd3_1
Xfanout904 net906 net904 VPWR VGND sg13g2_buf_8
Xfanout915 net917 net915 VPWR VGND sg13g2_buf_8
XFILLER_97_261 VPWR VGND sg13g2_decap_8
Xfanout948 net949 net948 VPWR VGND sg13g2_buf_8
Xfanout937 net938 net937 VPWR VGND sg13g2_buf_8
Xfanout926 net928 net926 VPWR VGND sg13g2_buf_8
Xhold1124 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[21\]
+ VPWR VGND net2951 sg13g2_dlygate4sd3_1
X_08824_ net1584 VGND VPWR _00882_ i_exotiny.i_wb_spi.state_r\[23\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
Xhold1102 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[8\]
+ VPWR VGND net2929 sg13g2_dlygate4sd3_1
Xfanout959 net960 net959 VPWR VGND sg13g2_buf_2
Xhold1113 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[19\]
+ VPWR VGND net2940 sg13g2_dlygate4sd3_1
XFILLER_38_28 VPWR VGND sg13g2_fill_1
X_08755_ net1653 VGND VPWR net3046 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[18\]
+ clknet_leaf_85_clk_regs sg13g2_dfrbpq_1
Xhold1157 _00559_ VPWR VGND net2984 sg13g2_dlygate4sd3_1
Xhold1146 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[26\]
+ VPWR VGND net2973 sg13g2_dlygate4sd3_1
Xhold1135 _00284_ VPWR VGND net2962 sg13g2_dlygate4sd3_1
XFILLER_94_990 VPWR VGND sg13g2_decap_8
Xhold1168 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[24\]
+ VPWR VGND net2995 sg13g2_dlygate4sd3_1
X_05967_ i_exotiny._0020_\[2\] net878 _02486_ _02490_ VPWR VGND sg13g2_mux2_1
XFILLER_72_106 VPWR VGND sg13g2_fill_2
X_07706_ net3490 net3459 net996 _01202_ VPWR VGND sg13g2_mux2_1
Xhold1179 i_exotiny._0024_\[1\] VPWR VGND net3006 sg13g2_dlygate4sd3_1
X_07899__45 VPWR VGND net45 sg13g2_tiehi
X_05898_ i_exotiny._0019_\[3\] net2895 net977 _00115_ VPWR VGND sg13g2_mux2_1
X_04918_ net1255 _01620_ _01640_ _01650_ VPWR VGND sg13g2_nor3_2
X_08686_ net1722 VGND VPWR net2989 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[13\]
+ clknet_leaf_116_clk_regs sg13g2_dfrbpq_1
X_04849_ _01572_ _01586_ _01587_ VPWR VGND sg13g2_nor2b_1
XFILLER_53_375 VPWR VGND sg13g2_fill_1
XFILLER_53_353 VPWR VGND sg13g2_fill_1
X_07637_ net2686 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[14\]
+ net897 _01145_ VPWR VGND sg13g2_mux2_1
XFILLER_41_515 VPWR VGND sg13g2_decap_4
X_07568_ i_exotiny._1737_ _01527_ _01545_ _03150_ _03151_ VPWR VGND sg13g2_nor4_1
XFILLER_13_217 VPWR VGND sg13g2_fill_1
X_06519_ net3153 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[12\]
+ net932 _00594_ VPWR VGND sg13g2_mux2_1
XFILLER_103_1007 VPWR VGND sg13g2_decap_8
XFILLER_10_935 VPWR VGND sg13g2_decap_8
X_07499_ net3661 net3665 net902 _01082_ VPWR VGND sg13g2_mux2_1
XFILLER_6_906 VPWR VGND sg13g2_decap_8
X_09238_ net699 VGND VPWR net3018 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[28\]
+ clknet_leaf_135_clk_regs sg13g2_dfrbpq_1
X_09169_ net813 VGND VPWR net2380 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[25\]
+ clknet_leaf_174_clk_regs sg13g2_dfrbpq_1
Xclkbuf_leaf_77_clk_regs clknet_5_26__leaf_clk_regs clknet_leaf_77_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold980 _00820_ VPWR VGND net2807 sg13g2_dlygate4sd3_1
Xhold991 _00122_ VPWR VGND net2818 sg13g2_dlygate4sd3_1
XFILLER_88_261 VPWR VGND sg13g2_fill_2
XFILLER_103_594 VPWR VGND sg13g2_fill_1
XFILLER_95_34 VPWR VGND sg13g2_fill_1
XFILLER_89_795 VPWR VGND sg13g2_fill_1
XFILLER_0_165 VPWR VGND sg13g2_fill_1
XFILLER_92_949 VPWR VGND sg13g2_decap_8
Xhold1680 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[30\]
+ VPWR VGND net3507 sg13g2_dlygate4sd3_1
XFILLER_29_350 VPWR VGND sg13g2_fill_2
XFILLER_56_191 VPWR VGND sg13g2_fill_2
XFILLER_17_523 VPWR VGND sg13g2_fill_1
Xhold1691 _00635_ VPWR VGND net3518 sg13g2_dlygate4sd3_1
XFILLER_72_684 VPWR VGND sg13g2_fill_2
X_08778__1210 VPWR VGND net1630 sg13g2_tiehi
X_08701__1287 VPWR VGND net1707 sg13g2_tiehi
XFILLER_5_994 VPWR VGND sg13g2_decap_8
X_06870_ net1172 VPWR _02879_ VGND net3623 net1186 sg13g2_o21ai_1
XFILLER_39_103 VPWR VGND sg13g2_fill_1
X_05821_ net2745 net2750 net1056 _00093_ VPWR VGND sg13g2_mux2_1
X_05752_ _02386_ net3636 _02384_ VPWR VGND sg13g2_xnor2_1
X_08923__1059 VPWR VGND net1479 sg13g2_tiehi
X_08540_ net140 VGND VPWR _00614_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[28\]
+ clknet_leaf_177_clk_regs sg13g2_dfrbpq_1
X_05683_ net1926 net1063 _02333_ VPWR VGND sg13g2_nor2_1
X_08471_ net209 VGND VPWR net3116 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[23\]
+ clknet_leaf_158_clk_regs sg13g2_dfrbpq_1
X_04703_ net1253 _01460_ _01461_ VPWR VGND sg13g2_nor2b_2
X_04634_ VPWR _01396_ net3838 VGND sg13g2_inv_1
X_07422_ net1083 _03067_ _03068_ _03069_ VPWR VGND sg13g2_nor3_1
XFILLER_50_389 VPWR VGND sg13g2_fill_2
X_07353_ _03015_ _03004_ net2997 VPWR VGND sg13g2_nand2b_1
X_07284_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[9\]
+ net2067 net908 _01001_ VPWR VGND sg13g2_mux2_1
X_06304_ _02420_ _02525_ _02558_ VPWR VGND sg13g2_nor2_2
X_06235_ net2416 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[5\]
+ net1040 _00384_ VPWR VGND sg13g2_mux2_1
X_09023_ net1379 VGND VPWR _01081_ i_exotiny._0315_\[11\] clknet_leaf_179_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_105_804 VPWR VGND sg13g2_decap_8
XFILLER_85_1013 VPWR VGND sg13g2_decap_8
Xhold210 i_exotiny._0314_\[31\] VPWR VGND net2037 sg13g2_dlygate4sd3_1
X_06166_ net3149 net3441 net952 _00328_ VPWR VGND sg13g2_mux2_1
Xhold243 _01329_ VPWR VGND net2070 sg13g2_dlygate4sd3_1
Xhold221 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[24\]
+ VPWR VGND net2048 sg13g2_dlygate4sd3_1
Xhold232 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[4\]
+ VPWR VGND net2059 sg13g2_dlygate4sd3_1
Xhold276 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[25\]
+ VPWR VGND net2103 sg13g2_dlygate4sd3_1
Xhold265 _00107_ VPWR VGND net2092 sg13g2_dlygate4sd3_1
X_06097_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[23\]
+ net2435 net958 _00273_ VPWR VGND sg13g2_mux2_1
Xhold254 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[7\]
+ VPWR VGND net2081 sg13g2_dlygate4sd3_1
Xhold287 _00460_ VPWR VGND net2114 sg13g2_dlygate4sd3_1
X_05117_ _01847_ i_exotiny._0032_\[2\] _01767_ VPWR VGND sg13g2_nand2_1
XFILLER_104_369 VPWR VGND sg13g2_decap_8
Xhold298 i_exotiny._0369_\[21\] VPWR VGND net2125 sg13g2_dlygate4sd3_1
X_05048_ net1236 _01753_ _01757_ _01780_ VPWR VGND sg13g2_nor3_2
XFILLER_59_957 VPWR VGND sg13g2_fill_1
X_08807_ net1601 VGND VPWR _00865_ i_exotiny.i_wb_spi.state_r\[6\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
X_09140__842 VPWR VGND net842 sg13g2_tiehi
X_06999_ i_exotiny._0032_\[3\] net2093 net918 _00766_ VPWR VGND sg13g2_mux2_1
X_08738_ net1670 VGND VPWR _00796_ i_exotiny._0017_\[1\] clknet_leaf_81_clk_regs sg13g2_dfrbpq_2
XFILLER_85_297 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_124_clk_regs clknet_5_23__leaf_clk_regs clknet_leaf_124_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_38_191 VPWR VGND sg13g2_fill_1
XFILLER_45_128 VPWR VGND sg13g2_fill_1
X_08669_ net1203 VGND VPWR i_exotiny._2043_\[6\] i_exotiny._2034_\[6\] net1229 sg13g2_dfrbpq_2
XFILLER_92_1028 VPWR VGND sg13g2_fill_1
XFILLER_14_96 VPWR VGND sg13g2_fill_2
XFILLER_22_592 VPWR VGND sg13g2_fill_2
XFILLER_10_798 VPWR VGND sg13g2_decap_4
XFILLER_30_40 VPWR VGND sg13g2_fill_1
XFILLER_100_0 VPWR VGND sg13g2_fill_2
XFILLER_5_268 VPWR VGND sg13g2_fill_1
XFILLER_96_507 VPWR VGND sg13g2_decap_8
XFILLER_1_430 VPWR VGND sg13g2_fill_1
XFILLER_2_964 VPWR VGND sg13g2_decap_8
XFILLER_104_881 VPWR VGND sg13g2_decap_8
XFILLER_7_1024 VPWR VGND sg13g2_decap_4
XFILLER_1_485 VPWR VGND sg13g2_fill_2
XFILLER_39_82 VPWR VGND sg13g2_decap_8
XFILLER_36_139 VPWR VGND sg13g2_fill_1
X_08719__1269 VPWR VGND net1689 sg13g2_tiehi
XFILLER_13_570 VPWR VGND sg13g2_fill_2
XFILLER_32_367 VPWR VGND sg13g2_fill_1
XFILLER_9_596 VPWR VGND sg13g2_fill_1
X_06020_ VGND VPWR net3559 net1103 _00212_ _02504_ sg13g2_a21oi_1
XFILLER_102_818 VPWR VGND sg13g2_decap_8
XFILLER_99_367 VPWR VGND sg13g2_decap_8
X_07971_ net1177 VGND VPWR net1876 i_exotiny.i_wdg_top.o_wb_dat\[12\] clknet_leaf_57_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_101_317 VPWR VGND sg13g2_decap_8
X_06922_ i_exotiny._0029_\[2\] net2408 net926 _00701_ VPWR VGND sg13g2_mux2_1
X_06853_ net1129 _02863_ _02864_ _02865_ VPWR VGND sg13g2_nor3_1
XFILLER_55_415 VPWR VGND sg13g2_fill_2
X_06784_ net1171 VPWR _02807_ VGND net1945 _01451_ sg13g2_o21ai_1
XFILLER_55_448 VPWR VGND sg13g2_fill_2
X_05804_ _02419_ _02420_ _02421_ VPWR VGND sg13g2_nor2_2
X_05735_ _02372_ i_exotiny.i_wb_regs.spi_size_o\[0\] i_exotiny.i_wb_regs.spi_size_o\[1\]
+ VPWR VGND sg13g2_nand2_1
X_08523_ net157 VGND VPWR _00597_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[11\]
+ clknet_leaf_182_clk_regs sg13g2_dfrbpq_1
X_08662__775 VPWR VGND net775 sg13g2_tiehi
X_05666_ VGND VPWR net1064 _02319_ _00042_ _02320_ sg13g2_a21oi_1
X_08454_ net226 VGND VPWR _00528_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[6\]
+ clknet_leaf_114_clk_regs sg13g2_dfrbpq_1
XFILLER_50_120 VPWR VGND sg13g2_fill_1
X_04617_ VPWR _01379_ net3634 VGND sg13g2_inv_1
XFILLER_51_676 VPWR VGND sg13g2_fill_2
X_07405_ VGND VPWR i_exotiny._0369_\[13\] net1147 _03056_ _03052_ sg13g2_a21oi_1
X_08385_ net293 VGND VPWR _00466_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[23\]
+ clknet_leaf_140_clk_regs sg13g2_dfrbpq_1
X_05597_ _01473_ _02260_ ccx_req VPWR VGND sg13g2_nor2_1
X_07336_ _03000_ i_exotiny._0369_\[6\] _02994_ VPWR VGND sg13g2_nand2_1
XFILLER_13_1018 VPWR VGND sg13g2_decap_8
X_07267_ i_exotiny._0040_\[1\] net883 _02972_ _02975_ VPWR VGND sg13g2_mux2_1
X_09006_ net1396 VGND VPWR net1912 i_exotiny._1160_\[27\] clknet_leaf_14_clk_regs
+ sg13g2_dfrbpq_1
X_07198_ net1967 net1092 _02961_ VPWR VGND sg13g2_nor2_1
X_06218_ net2671 net2774 net945 _00373_ VPWR VGND sg13g2_mux2_1
X_06149_ _02532_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[3\] i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[4\]
+ VPWR VGND sg13g2_nand2_2
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_105_678 VPWR VGND sg13g2_decap_8
XFILLER_104_166 VPWR VGND sg13g2_decap_8
XFILLER_74_713 VPWR VGND sg13g2_fill_2
XFILLER_18_128 VPWR VGND sg13g2_fill_2
XFILLER_92_68 VPWR VGND sg13g2_fill_2
XFILLER_70_974 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_92_clk_regs clknet_5_31__leaf_clk_regs clknet_leaf_92_clk_regs VPWR VGND
+ sg13g2_buf_8
Xclkbuf_leaf_21_clk_regs clknet_5_12__leaf_clk_regs clknet_leaf_21_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_97_805 VPWR VGND sg13g2_fill_2
XFILLER_97_849 VPWR VGND sg13g2_decap_8
XFILLER_96_315 VPWR VGND sg13g2_decap_8
XFILLER_69_529 VPWR VGND sg13g2_fill_2
XFILLER_2_761 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_17_161 VPWR VGND sg13g2_fill_1
XFILLER_61_974 VPWR VGND sg13g2_fill_1
X_05520_ net1275 i_exotiny._0315_\[13\] _02210_ VPWR VGND sg13g2_nor2b_1
X_05451_ VPWR VGND i_exotiny._1617_\[1\] _02158_ _02149_ i_exotiny._1612_\[1\] _02159_
+ _02148_ sg13g2_a221oi_1
XFILLER_33_676 VPWR VGND sg13g2_fill_2
X_08170_ net507 VGND VPWR _00251_ i_exotiny._0038_\[1\] clknet_leaf_112_clk_regs sg13g2_dfrbpq_2
X_08855__1131 VPWR VGND net1551 sg13g2_tiehi
X_07121_ net1290 net1849 _00871_ VPWR VGND sg13g2_and2_1
X_05382_ _02093_ net1112 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set[0]
+ _02103_ VPWR VGND sg13g2_a21o_1
X_09130__852 VPWR VGND net852 sg13g2_tiehi
X_07052_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[22\]
+ net3045 net1017 _00813_ VPWR VGND sg13g2_mux2_1
X_06003_ net3513 _02495_ net1049 _00204_ VPWR VGND sg13g2_mux2_1
X_07954_ net1179 VGND VPWR i_exotiny._2055_\[2\] i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_hw_set[0]
+ clknet_leaf_40_clk_regs sg13g2_dfrbpq_2
XFILLER_96_893 VPWR VGND sg13g2_decap_8
X_06905_ _02905_ _02903_ net1227 _02906_ VPWR VGND sg13g2_a21o_1
X_07885_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[23\]
+ net2190 _03229_ _01352_ VPWR VGND sg13g2_mux2_1
X_07992__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_28_404 VPWR VGND sg13g2_fill_1
XFILLER_95_392 VPWR VGND sg13g2_decap_4
X_06836_ VGND VPWR i_exotiny._1616_\[2\] net1132 _02851_ _02850_ sg13g2_a21oi_1
X_07944__88 VPWR VGND net88 sg13g2_tiehi
XFILLER_55_267 VPWR VGND sg13g2_fill_2
X_06767_ net2331 net1100 _02793_ VPWR VGND sg13g2_nor2_1
XFILLER_83_587 VPWR VGND sg13g2_fill_1
XFILLER_55_278 VPWR VGND sg13g2_fill_2
X_08506_ net174 VGND VPWR _00580_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[26\]
+ clknet_leaf_71_clk_regs sg13g2_dfrbpq_1
XFILLER_70_248 VPWR VGND sg13g2_fill_2
X_05718_ VGND VPWR net1059 _02359_ _00055_ _02357_ sg13g2_a21oi_1
X_06698_ _02734_ _02723_ net16 _02593_ net3618 VPWR VGND sg13g2_a22oi_1
X_08660__1317 VPWR VGND net1737 sg13g2_tiehi
XFILLER_36_492 VPWR VGND sg13g2_fill_1
X_05649_ net1953 net1066 _02308_ VPWR VGND sg13g2_nor2_1
X_08437_ net248 VGND VPWR _00511_ i_exotiny._0369_\[8\] clknet_leaf_16_clk_regs sg13g2_dfrbpq_2
XFILLER_23_175 VPWR VGND sg13g2_fill_1
XFILLER_11_359 VPWR VGND sg13g2_fill_2
X_08368_ net310 VGND VPWR _00449_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[6\]
+ clknet_leaf_137_clk_regs sg13g2_dfrbpq_1
X_08299_ net379 VGND VPWR net3516 i_exotiny._0031_\[1\] clknet_leaf_72_clk_regs sg13g2_dfrbpq_2
X_08539__141 VPWR VGND net141 sg13g2_tiehi
X_07319_ _02986_ net3749 net1150 VPWR VGND sg13g2_nand2_1
XFILLER_106_965 VPWR VGND sg13g2_decap_8
XFILLER_105_431 VPWR VGND sg13g2_decap_8
XFILLER_79_805 VPWR VGND sg13g2_fill_1
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_4_1016 VPWR VGND sg13g2_decap_8
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
XFILLER_59_1007 VPWR VGND sg13g2_fill_1
XFILLER_62_738 VPWR VGND sg13g2_fill_1
XFILLER_61_248 VPWR VGND sg13g2_decap_4
X_08636__1341 VPWR VGND net1761 sg13g2_tiehi
XFILLER_43_985 VPWR VGND sg13g2_fill_2
XFILLER_30_646 VPWR VGND sg13g2_fill_1
Xinput14 uio_in[4] net14 VPWR VGND sg13g2_buf_2
X_09291__1397 VPWR VGND net1817 sg13g2_tiehi
XFILLER_7_886 VPWR VGND sg13g2_fill_2
Xhold809 _00699_ VPWR VGND net2636 sg13g2_dlygate4sd3_1
X_07976__117 VPWR VGND net117 sg13g2_tiehi
XFILLER_35_4 VPWR VGND sg13g2_fill_1
Xhold1509 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[6\]
+ VPWR VGND net3336 sg13g2_dlygate4sd3_1
X_04951_ _01683_ _01427_ _01429_ VPWR VGND sg13g2_nand2_1
X_04882_ i_exotiny._0077_\[2\] i_exotiny._0077_\[3\] net1223 _01614_ VPWR VGND sg13g2_or3_1
X_07670_ net2535 net2301 net998 _01172_ VPWR VGND sg13g2_mux2_1
X_06621_ net1198 _02669_ _02670_ _00647_ VPWR VGND sg13g2_nor3_1
X_06552_ net3443 net1213 _02628_ VPWR VGND sg13g2_and2_1
X_05503_ _02197_ net3505 net1069 VPWR VGND sg13g2_nand2_1
X_09271_ net79 VGND VPWR net2911 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[29\]
+ clknet_leaf_127_clk_regs sg13g2_dfrbpq_1
X_06483_ net3298 net2530 net1026 _00564_ VPWR VGND sg13g2_mux2_1
XFILLER_60_270 VPWR VGND sg13g2_fill_2
X_08222_ net455 VGND VPWR _00303_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[21\]
+ clknet_leaf_153_clk_regs sg13g2_dfrbpq_1
X_05434_ VPWR _02143_ _02142_ VGND sg13g2_inv_1
X_05365_ VGND VPWR _00014_ i_exotiny._2034_\[0\] _02087_ _02080_ sg13g2_a21oi_1
X_08153_ net525 VGND VPWR _00234_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[17\]
+ clknet_leaf_133_clk_regs sg13g2_dfrbpq_1
X_08084_ net610 VGND VPWR net2459 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[21\]
+ clknet_leaf_92_clk_regs sg13g2_dfrbpq_1
X_07104_ net3080 net876 _02940_ _02944_ VPWR VGND sg13g2_mux2_1
X_07035_ net3593 net3129 net1014 _00796_ VPWR VGND sg13g2_mux2_1
X_05296_ _02022_ _01636_ i_exotiny._0019_\[0\] _01628_ i_exotiny._0037_\[0\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_103_902 VPWR VGND sg13g2_decap_8
X_08176__501 VPWR VGND net501 sg13g2_tiehi
XFILLER_0_517 VPWR VGND sg13g2_fill_2
XFILLER_102_434 VPWR VGND sg13g2_decap_8
X_08986_ net1416 VGND VPWR net1956 i_exotiny._1160_\[7\] clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
XFILLER_103_979 VPWR VGND sg13g2_decap_8
X_07937_ net711 VGND VPWR net1999 i_exotiny._1924_\[30\] clknet_leaf_30_clk_regs sg13g2_dfrbpq_1
XFILLER_57_49 VPWR VGND sg13g2_fill_2
X_08714__1274 VPWR VGND net1694 sg13g2_tiehi
X_07868_ net2451 net3268 net981 _01335_ VPWR VGND sg13g2_mux2_1
X_06819_ net3711 net1097 _02837_ VPWR VGND sg13g2_nor2_1
X_07799_ net3340 net2625 net894 _01278_ VPWR VGND sg13g2_mux2_1
XFILLER_25_963 VPWR VGND sg13g2_fill_1
X_08936__1046 VPWR VGND net1466 sg13g2_tiehi
XFILLER_7_105 VPWR VGND sg13g2_fill_2
XFILLER_4_834 VPWR VGND sg13g2_decap_8
X_08296__382 VPWR VGND net382 sg13g2_tiehi
XFILLER_106_762 VPWR VGND sg13g2_decap_8
Xfanout1112 _02091_ net1112 VPWR VGND sg13g2_buf_8
Xfanout1101 net1102 net1101 VPWR VGND sg13g2_buf_8
Xfanout1145 _01549_ net1145 VPWR VGND sg13g2_buf_8
Xfanout1123 _01582_ net1123 VPWR VGND sg13g2_buf_8
Xfanout1134 net1135 net1134 VPWR VGND sg13g2_buf_8
Xfanout1156 net1157 net1156 VPWR VGND sg13g2_buf_2
Xfanout1178 net1179 net1178 VPWR VGND sg13g2_buf_8
Xfanout1189 _01450_ net1189 VPWR VGND sg13g2_buf_2
Xfanout1167 net1168 net1167 VPWR VGND sg13g2_buf_1
X_09120__862 VPWR VGND net862 sg13g2_tiehi
X_08444__238 VPWR VGND net238 sg13g2_tiehi
X_05150_ _01880_ _01638_ i_exotiny._0029_\[2\] _01625_ i_exotiny._0030_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold606 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[23\]
+ VPWR VGND net2433 sg13g2_dlygate4sd3_1
Xhold617 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[29\]
+ VPWR VGND net2444 sg13g2_dlygate4sd3_1
Xhold628 _00979_ VPWR VGND net2455 sg13g2_dlygate4sd3_1
Xhold639 _00444_ VPWR VGND net2466 sg13g2_dlygate4sd3_1
X_05081_ _01812_ VPWR _01813_ VGND i_exotiny._0036_\[3\] _01755_ sg13g2_o21ai_1
XFILLER_98_944 VPWR VGND sg13g2_decap_8
XFILLER_97_443 VPWR VGND sg13g2_decap_8
X_08840_ net1566 VGND VPWR _00898_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[7\]
+ clknet_leaf_185_clk_regs sg13g2_dfrbpq_1
Xhold2007 i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[2\] VPWR VGND net3834 sg13g2_dlygate4sd3_1
Xhold1306 i_exotiny._0041_\[1\] VPWR VGND net3133 sg13g2_dlygate4sd3_1
XFILLER_26_0 VPWR VGND sg13g2_decap_4
XFILLER_100_938 VPWR VGND sg13g2_decap_8
Xhold1317 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[2\] VPWR VGND net3144
+ sg13g2_dlygate4sd3_1
X_05983_ net2586 net2595 net1050 _00185_ VPWR VGND sg13g2_mux2_1
Xhold1328 i_exotiny._0314_\[23\] VPWR VGND net3155 sg13g2_dlygate4sd3_1
X_08771_ net1637 VGND VPWR _00829_ i_exotiny._0015_\[2\] clknet_leaf_158_clk_regs
+ sg13g2_dfrbpq_2
Xhold1339 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[23\]
+ VPWR VGND net3166 sg13g2_dlygate4sd3_1
XFILLER_66_863 VPWR VGND sg13g2_fill_1
X_07722_ net2885 net2568 net995 _01218_ VPWR VGND sg13g2_mux2_1
X_04934_ VPWR VGND i_exotiny._0025_\[3\] _01665_ _01645_ i_exotiny._0023_\[3\] _01666_
+ _01622_ sg13g2_a221oi_1
X_07653_ net3004 net2296 net897 _01161_ VPWR VGND sg13g2_mux2_1
X_08529__151 VPWR VGND net151 sg13g2_tiehi
X_04865_ net1268 i_exotiny._1306_ _01598_ VPWR VGND sg13g2_nor2_2
XFILLER_38_598 VPWR VGND sg13g2_fill_1
X_06604_ i_exotiny._0314_\[14\] net1163 _02659_ VPWR VGND sg13g2_nor2_1
XFILLER_25_237 VPWR VGND sg13g2_fill_1
X_07584_ _03161_ net3671 _03159_ VPWR VGND sg13g2_xnor2_1
XFILLER_80_365 VPWR VGND sg13g2_fill_1
X_04796_ VGND VPWR _01543_ _01544_ _00011_ _01487_ sg13g2_a21oi_1
X_06535_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[24\]
+ net2617 net933 _00610_ VPWR VGND sg13g2_mux2_1
XFILLER_40_218 VPWR VGND sg13g2_fill_2
X_06466_ _02611_ net2249 net936 _00551_ VPWR VGND sg13g2_mux2_1
X_09254_ net553 VGND VPWR net2809 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[12\]
+ clknet_leaf_128_clk_regs sg13g2_dfrbpq_1
X_09185_ net796 VGND VPWR net2461 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[7\]
+ clknet_leaf_76_clk_regs sg13g2_dfrbpq_1
X_05417_ _01529_ VPWR _02126_ VGND i_exotiny._0327_\[0\] _01533_ sg13g2_o21ai_1
X_08205_ net472 VGND VPWR _00286_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[4\]
+ clknet_leaf_151_clk_regs sg13g2_dfrbpq_1
XFILLER_88_1000 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_149_clk_regs clknet_5_16__leaf_clk_regs clknet_leaf_149_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08136_ net549 VGND VPWR net2638 i_exotiny._0025_\[0\] clknet_leaf_120_clk_regs sg13g2_dfrbpq_2
X_06397_ _00511_ net1284 net3829 VPWR VGND sg13g2_nand2_1
X_05348_ i_exotiny.i_wb_regs.spi_auto_cs_o _02070_ _02071_ VPWR VGND i_exotiny.gpo\[1\]
+ sg13g2_nand3b_1
X_08067_ net627 VGND VPWR net2320 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[4\]
+ clknet_leaf_89_clk_regs sg13g2_dfrbpq_1
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
X_08536__144 VPWR VGND net144 sg13g2_tiehi
X_05279_ _02005_ _01780_ i_exotiny._0041_\[0\] _01763_ i_exotiny._0029_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_07018_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[22\]
+ net2111 net920 _00785_ VPWR VGND sg13g2_mux2_1
XFILLER_1_859 VPWR VGND sg13g2_decap_8
XFILLER_103_776 VPWR VGND sg13g2_decap_8
XFILLER_102_231 VPWR VGND sg13g2_decap_8
XFILLER_89_988 VPWR VGND sg13g2_decap_8
XFILLER_49_819 VPWR VGND sg13g2_fill_1
X_08969_ net1433 VGND VPWR _01027_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[5\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
Xhold1840 _00068_ VPWR VGND net3667 sg13g2_dlygate4sd3_1
Xhold1862 _02597_ VPWR VGND net3689 sg13g2_dlygate4sd3_1
Xhold1851 _02248_ VPWR VGND net3678 sg13g2_dlygate4sd3_1
Xhold1895 i_exotiny.i_wdg_top.clk_div_inst.cnt\[14\] VPWR VGND net3722 sg13g2_dlygate4sd3_1
Xhold1884 i_exotiny._1614_\[3\] VPWR VGND net3711 sg13g2_dlygate4sd3_1
Xhold1873 _03152_ VPWR VGND net3700 sg13g2_dlygate4sd3_1
XFILLER_8_447 VPWR VGND sg13g2_fill_1
XFILLER_79_465 VPWR VGND sg13g2_fill_2
Xhold3 i_exotiny.i_wdg_top.clk_div_inst.cnt\[0\] VPWR VGND net1830 sg13g2_dlygate4sd3_1
XFILLER_95_947 VPWR VGND sg13g2_decap_8
XFILLER_82_608 VPWR VGND sg13g2_fill_1
XFILLER_94_479 VPWR VGND sg13g2_fill_2
XFILLER_74_80 VPWR VGND sg13g2_fill_1
X_04650_ VPWR _01412_ net2105 VGND sg13g2_inv_1
X_06320_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[18\]
+ net3257 net1036 _00457_ VPWR VGND sg13g2_mux2_1
X_06251_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[25\]
+ net2373 net1040 _00400_ VPWR VGND sg13g2_mux2_1
X_05202_ _01925_ _01928_ _01923_ _01930_ VPWR VGND _01929_ sg13g2_nand4_1
X_06182_ net885 i_exotiny._0028_\[1\] _02533_ _02536_ VPWR VGND sg13g2_mux2_1
Xhold414 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[17\]
+ VPWR VGND net2241 sg13g2_dlygate4sd3_1
Xhold436 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[19\]
+ VPWR VGND net2263 sg13g2_dlygate4sd3_1
Xhold403 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[5\]
+ VPWR VGND net2230 sg13g2_dlygate4sd3_1
Xhold425 _01276_ VPWR VGND net2252 sg13g2_dlygate4sd3_1
X_05133_ _01863_ _01786_ i_exotiny._0017_\[2\] _01782_ i_exotiny._0037_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold447 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[7\]
+ VPWR VGND net2274 sg13g2_dlygate4sd3_1
Xhold458 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[5\]
+ VPWR VGND net2285 sg13g2_dlygate4sd3_1
Xhold469 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[30\]
+ VPWR VGND net2296 sg13g2_dlygate4sd3_1
X_05064_ _01796_ _01773_ i_exotiny._0019_\[3\] _01761_ i_exotiny._0015_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_08173__504 VPWR VGND net504 sg13g2_tiehi
Xfanout905 net906 net905 VPWR VGND sg13g2_buf_1
Xfanout916 net917 net916 VPWR VGND sg13g2_buf_8
Xfanout949 _02541_ net949 VPWR VGND sg13g2_buf_8
Xfanout938 _02609_ net938 VPWR VGND sg13g2_buf_8
Xfanout927 net928 net927 VPWR VGND sg13g2_buf_8
X_08823_ net1585 VGND VPWR _00881_ i_exotiny.i_wb_spi.state_r\[22\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
Xhold1103 _00483_ VPWR VGND net2930 sg13g2_dlygate4sd3_1
Xhold1114 _00573_ VPWR VGND net2941 sg13g2_dlygate4sd3_1
XFILLER_100_746 VPWR VGND sg13g2_fill_1
X_09203__778 VPWR VGND net778 sg13g2_tiehi
X_08754_ net1654 VGND VPWR net2223 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[17\]
+ clknet_leaf_87_clk_regs sg13g2_dfrbpq_1
X_05966_ net2772 _02489_ net966 _00173_ VPWR VGND sg13g2_mux2_1
Xhold1136 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[18\]
+ VPWR VGND net2963 sg13g2_dlygate4sd3_1
XFILLER_57_159 VPWR VGND sg13g2_fill_1
Xhold1158 i_exotiny._0029_\[0\] VPWR VGND net2985 sg13g2_dlygate4sd3_1
Xhold1125 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[19\]
+ VPWR VGND net2952 sg13g2_dlygate4sd3_1
Xhold1147 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[27\]
+ VPWR VGND net2974 sg13g2_dlygate4sd3_1
Xhold1169 _00499_ VPWR VGND net2996 sg13g2_dlygate4sd3_1
X_04917_ net1258 net1260 net1255 _01649_ VGND VPWR _01616_ sg13g2_nor4_2
X_07705_ net2724 net2613 net996 _01201_ VPWR VGND sg13g2_mux2_1
X_05897_ i_exotiny._0019_\[2\] net2867 net976 _00114_ VPWR VGND sg13g2_mux2_1
X_08685_ net1723 VGND VPWR net2723 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[12\]
+ clknet_leaf_102_clk_regs sg13g2_dfrbpq_1
X_04848_ net3814 VPWR _01586_ VGND net1840 net3728 sg13g2_o21ai_1
X_07636_ net2607 net3190 net898 _01144_ VPWR VGND sg13g2_mux2_1
X_08286__392 VPWR VGND net392 sg13g2_tiehi
X_07567_ _01493_ net3520 _03146_ _03150_ VPWR VGND sg13g2_a21o_1
XFILLER_41_527 VPWR VGND sg13g2_fill_2
X_04779_ _01529_ net1224 net1234 VPWR VGND sg13g2_nand2_1
X_06518_ net2274 net2590 net930 _00593_ VPWR VGND sg13g2_mux2_1
X_07498_ net3612 net3626 net904 _01081_ VPWR VGND sg13g2_mux2_1
XFILLER_16_1027 VPWR VGND sg13g2_fill_2
XFILLER_21_240 VPWR VGND sg13g2_fill_2
X_09237_ net701 VGND VPWR net2498 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[27\]
+ clknet_leaf_133_clk_regs sg13g2_dfrbpq_1
X_06449_ net2648 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[14\]
+ net938 _00536_ VPWR VGND sg13g2_mux2_1
X_09168_ net814 VGND VPWR _01223_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[24\]
+ clknet_leaf_174_clk_regs sg13g2_dfrbpq_1
X_08119_ net575 VGND VPWR net2755 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[24\]
+ clknet_leaf_101_clk_regs sg13g2_dfrbpq_1
X_09110__872 VPWR VGND net1292 sg13g2_tiehi
X_09099_ net1303 VGND VPWR _01154_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[19\]
+ clknet_leaf_145_clk_regs sg13g2_dfrbpq_1
XFILLER_102_4 VPWR VGND sg13g2_fill_2
Xhold970 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[17\]
+ VPWR VGND net2797 sg13g2_dlygate4sd3_1
Xhold981 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[12\]
+ VPWR VGND net2808 sg13g2_dlygate4sd3_1
X_08886__1096 VPWR VGND net1516 sg13g2_tiehi
X_08293__385 VPWR VGND net385 sg13g2_tiehi
Xhold992 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[22\]
+ VPWR VGND net2819 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_46_clk_regs clknet_5_11__leaf_clk_regs clknet_leaf_46_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_76_468 VPWR VGND sg13g2_fill_1
XFILLER_92_928 VPWR VGND sg13g2_decap_8
Xhold1670 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[5\]
+ VPWR VGND net3497 sg13g2_dlygate4sd3_1
Xhold1692 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[6\]
+ VPWR VGND net3519 sg13g2_dlygate4sd3_1
Xhold1681 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[7\]
+ VPWR VGND net3508 sg13g2_dlygate4sd3_1
XFILLER_32_538 VPWR VGND sg13g2_fill_2
XFILLER_40_560 VPWR VGND sg13g2_decap_4
X_08673__1315 VPWR VGND net1735 sg13g2_tiehi
XFILLER_5_11 VPWR VGND sg13g2_decap_8
X_08519__161 VPWR VGND net161 sg13g2_tiehi
XFILLER_5_973 VPWR VGND sg13g2_decap_8
XFILLER_68_903 VPWR VGND sg13g2_fill_1
XFILLER_95_744 VPWR VGND sg13g2_fill_1
X_05820_ net2152 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[12\]
+ net1053 _00092_ VPWR VGND sg13g2_mux2_1
XFILLER_82_405 VPWR VGND sg13g2_fill_1
XFILLER_94_298 VPWR VGND sg13g2_decap_8
X_05751_ i_exotiny._1956_ i_exotiny.i_wb_spi.cnt_hbit_r\[1\] net1072 _02385_ VPWR
+ VGND sg13g2_nor3_1
X_08931__1051 VPWR VGND net1471 sg13g2_tiehi
X_05682_ VGND VPWR net1063 _02332_ _00046_ _02330_ sg13g2_a21oi_1
XFILLER_62_151 VPWR VGND sg13g2_fill_1
X_08470_ net210 VGND VPWR _00544_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[22\]
+ clknet_leaf_114_clk_regs sg13g2_dfrbpq_1
X_04702_ _01458_ net1242 _01459_ _01460_ VPWR VGND sg13g2_a21o_1
XFILLER_91_994 VPWR VGND sg13g2_decap_8
X_08526__154 VPWR VGND net154 sg13g2_tiehi
X_07421_ VGND VPWR i_exotiny._0369_\[17\] net1147 _03068_ _03052_ sg13g2_a21oi_1
X_04633_ VPWR _01395_ net1237 VGND sg13g2_inv_1
X_07352_ i_exotiny._0369_\[3\] _02998_ _03014_ VPWR VGND sg13g2_nor2_2
X_06303_ _02557_ net2673 net942 _00442_ VPWR VGND sg13g2_mux2_1
X_07283_ net2767 net3363 net910 _01000_ VPWR VGND sg13g2_mux2_1
X_06234_ net2986 net2095 net1040 _00383_ VPWR VGND sg13g2_mux2_1
X_09022_ net1380 VGND VPWR _01080_ i_exotiny._0315_\[10\] clknet_leaf_166_clk_regs
+ sg13g2_dfrbpq_1
X_06165_ net2218 net2873 net952 _00327_ VPWR VGND sg13g2_mux2_1
Xhold211 i_exotiny._0314_\[24\] VPWR VGND net2038 sg13g2_dlygate4sd3_1
Xhold200 _01043_ VPWR VGND net2027 sg13g2_dlygate4sd3_1
Xhold222 _01219_ VPWR VGND net2049 sg13g2_dlygate4sd3_1
Xhold244 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[8\]
+ VPWR VGND net2071 sg13g2_dlygate4sd3_1
X_05116_ i_exotiny._0036_\[2\] _01755_ _01846_ VPWR VGND sg13g2_nor2_1
Xhold233 _00763_ VPWR VGND net2060 sg13g2_dlygate4sd3_1
Xhold277 _01013_ VPWR VGND net2104 sg13g2_dlygate4sd3_1
X_06096_ net2413 net2769 net958 _00272_ VPWR VGND sg13g2_mux2_1
Xhold255 _00557_ VPWR VGND net2082 sg13g2_dlygate4sd3_1
X_08533__147 VPWR VGND net147 sg13g2_tiehi
Xhold266 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[7\]
+ VPWR VGND net2093 sg13g2_dlygate4sd3_1
XFILLER_104_348 VPWR VGND sg13g2_decap_8
XFILLER_59_914 VPWR VGND sg13g2_fill_2
Xhold288 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[7\]
+ VPWR VGND net2115 sg13g2_dlygate4sd3_1
Xhold299 i_exotiny._1611_\[17\] VPWR VGND net2126 sg13g2_dlygate4sd3_1
X_05047_ _01762_ _01768_ _01779_ VPWR VGND sg13g2_nor2_2
XFILLER_105_34 VPWR VGND sg13g2_fill_1
XFILLER_100_554 VPWR VGND sg13g2_fill_1
XFILLER_100_521 VPWR VGND sg13g2_decap_8
X_08806_ net1602 VGND VPWR _00864_ i_exotiny.i_wb_spi.state_r\[5\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_86_788 VPWR VGND sg13g2_fill_2
XFILLER_73_427 VPWR VGND sg13g2_fill_1
X_06998_ i_exotiny._0032_\[2\] net2627 net919 _00765_ VPWR VGND sg13g2_mux2_1
X_08737_ net1671 VGND VPWR net2411 i_exotiny._0017_\[0\] clknet_leaf_80_clk_regs sg13g2_dfrbpq_2
X_05949_ net2969 net3122 net967 _00158_ VPWR VGND sg13g2_mux2_1
X_08668_ i_exotiny.i_wdg_top.cntr_inst.rst_n_sync VGND VPWR i_exotiny._2043_\[5\]
+ i_exotiny._2034_\[5\] net1229 sg13g2_dfrbpq_2
X_08751__1237 VPWR VGND net1657 sg13g2_tiehi
X_07619_ net3569 _03182_ _03183_ VPWR VGND sg13g2_and2_1
X_08599_ net1797 VGND VPWR _00671_ i_exotiny._1612_\[3\] clknet_leaf_58_clk_regs sg13g2_dfrbpq_2
Xclkbuf_leaf_164_clk_regs clknet_5_4__leaf_clk_regs clknet_leaf_164_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08973__1009 VPWR VGND net1429 sg13g2_tiehi
XFILLER_2_943 VPWR VGND sg13g2_decap_8
XFILLER_30_96 VPWR VGND sg13g2_fill_1
XFILLER_104_860 VPWR VGND sg13g2_decap_8
XFILLER_77_733 VPWR VGND sg13g2_fill_2
XFILLER_7_1003 VPWR VGND sg13g2_decap_8
XFILLER_103_381 VPWR VGND sg13g2_decap_8
XFILLER_49_435 VPWR VGND sg13g2_fill_1
X_08727__1261 VPWR VGND net1681 sg13g2_tiehi
XFILLER_60_666 VPWR VGND sg13g2_fill_1
X_08622__1354 VPWR VGND net1774 sg13g2_tiehi
X_08949__1033 VPWR VGND net1453 sg13g2_tiehi
XFILLER_99_346 VPWR VGND sg13g2_decap_8
X_07970_ net1177 VGND VPWR net1871 i_exotiny.i_wdg_top.o_wb_dat\[11\] clknet_leaf_57_clk_regs
+ sg13g2_dfrbpq_1
X_06921_ i_exotiny._0029_\[1\] net2524 net924 _00700_ VPWR VGND sg13g2_mux2_1
X_08170__507 VPWR VGND net507 sg13g2_tiehi
XFILLER_56_917 VPWR VGND sg13g2_fill_1
X_06852_ net1170 VPWR _02864_ VGND i_exotiny.i_wb_spi.dat_rx_r\[25\] net1186 sg13g2_o21ai_1
X_06783_ net3643 net1191 _02806_ VPWR VGND sg13g2_nor2_1
X_05803_ _02420_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[3\] VPWR VGND
+ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[4\] sg13g2_nand2b_2
X_05734_ _02369_ VPWR _00059_ VGND net1073 _02371_ sg13g2_o21ai_1
X_08522_ net158 VGND VPWR _00596_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[10\]
+ clknet_leaf_183_clk_regs sg13g2_dfrbpq_1
X_09100__882 VPWR VGND net1302 sg13g2_tiehi
X_08453_ net227 VGND VPWR _00527_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[5\]
+ clknet_leaf_159_clk_regs sg13g2_dfrbpq_1
X_05665_ net2031 net1064 _02320_ VPWR VGND sg13g2_nor2_1
X_07404_ net2010 net1216 _03055_ VPWR VGND sg13g2_nor2_1
X_04616_ VPWR _01378_ net1291 VGND sg13g2_inv_1
X_08384_ net294 VGND VPWR net2017 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[22\]
+ clknet_leaf_134_clk_regs sg13g2_dfrbpq_1
X_05596_ _01834_ VPWR i_exotiny._1206_ VGND _01837_ _02268_ sg13g2_o21ai_1
X_08283__395 VPWR VGND net395 sg13g2_tiehi
Xclkbuf_0_clk_regs clk_regs clknet_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_50_176 VPWR VGND sg13g2_fill_1
X_07335_ _02999_ _02997_ _02998_ VPWR VGND sg13g2_nand2_2
X_07266_ _02974_ net3071 net1007 _00988_ VPWR VGND sg13g2_mux2_1
X_06217_ net2305 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[25\]
+ net945 _00372_ VPWR VGND sg13g2_mux2_1
X_09005_ net1397 VGND VPWR net3416 i_exotiny._1160_\[26\] clknet_leaf_165_clk_regs
+ sg13g2_dfrbpq_1
X_07197_ net3654 net1967 net1093 _00933_ VPWR VGND sg13g2_mux2_1
X_06148_ _02531_ net2658 net1046 _00313_ VPWR VGND sg13g2_mux2_1
XFILLER_105_657 VPWR VGND sg13g2_decap_8
XFILLER_104_145 VPWR VGND sg13g2_decap_8
X_06079_ net3091 net3193 net955 _00255_ VPWR VGND sg13g2_mux2_1
X_08769__1219 VPWR VGND net1639 sg13g2_tiehi
X_08805__1183 VPWR VGND net1603 sg13g2_tiehi
XFILLER_99_891 VPWR VGND sg13g2_decap_8
XFILLER_98_390 VPWR VGND sg13g2_decap_8
X_08290__388 VPWR VGND net388 sg13g2_tiehi
XFILLER_101_885 VPWR VGND sg13g2_decap_8
XFILLER_100_395 VPWR VGND sg13g2_decap_8
X_08509__171 VPWR VGND net171 sg13g2_tiehi
XFILLER_54_460 VPWR VGND sg13g2_decap_4
XFILLER_26_173 VPWR VGND sg13g2_fill_2
XFILLER_10_596 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_61_clk_regs clknet_5_13__leaf_clk_regs clknet_leaf_61_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08516__164 VPWR VGND net164 sg13g2_tiehi
XFILLER_49_232 VPWR VGND sg13g2_fill_2
XFILLER_77_596 VPWR VGND sg13g2_fill_2
XFILLER_64_213 VPWR VGND sg13g2_fill_1
X_05450_ _02156_ _02157_ _02155_ _02158_ VPWR VGND sg13g2_nand3_1
X_08523__157 VPWR VGND net157 sg13g2_tiehi
XFILLER_21_828 VPWR VGND sg13g2_fill_1
X_05381_ i_exotiny._2055_\[0\] _02100_ _02102_ _02073_ net3781 VPWR VGND sg13g2_a22oi_1
X_07120_ net1288 net1858 _00870_ VPWR VGND sg13g2_and2_1
XFILLER_9_383 VPWR VGND sg13g2_fill_1
X_07051_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[21\]
+ net2222 net1015 _00812_ VPWR VGND sg13g2_mux2_1
X_06002_ i_exotiny._0013_\[0\] net887 _02493_ _02495_ VPWR VGND sg13g2_mux2_1
XFILLER_88_828 VPWR VGND sg13g2_fill_1
XFILLER_87_327 VPWR VGND sg13g2_fill_1
X_08098__596 VPWR VGND net596 sg13g2_tiehi
X_07953_ net1179 VGND VPWR net1833 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_hw_set[0]
+ clknet_leaf_40_clk_regs sg13g2_dfrbpq_1
XFILLER_96_872 VPWR VGND sg13g2_decap_8
X_06904_ net2570 net1883 _01389_ _02904_ _02905_ VPWR VGND sg13g2_nor4_1
XFILLER_83_500 VPWR VGND sg13g2_decap_4
X_07884_ net2259 net3150 net982 _01351_ VPWR VGND sg13g2_mux2_1
XFILLER_95_382 VPWR VGND sg13g2_decap_4
X_06835_ net1129 _02848_ _02849_ _02850_ VPWR VGND sg13g2_nor3_1
X_06766_ VGND VPWR net3801 net1135 _02792_ _02791_ sg13g2_a21oi_1
X_08505_ net175 VGND VPWR _00579_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[25\]
+ clknet_leaf_71_clk_regs sg13g2_dfrbpq_1
X_05717_ VGND VPWR i_exotiny._1618_\[1\] net1114 _02359_ _02358_ sg13g2_a21oi_1
X_06697_ _02733_ net3576 net1193 VPWR VGND sg13g2_nand2_1
X_05648_ VGND VPWR i_exotiny._1614_\[0\] net1125 _02307_ _02306_ sg13g2_a21oi_1
XFILLER_24_688 VPWR VGND sg13g2_fill_2
X_08436_ net249 VGND VPWR _00510_ i_exotiny._0369_\[20\] clknet_leaf_15_clk_regs sg13g2_dfrbpq_2
X_08367_ net311 VGND VPWR _00448_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[5\]
+ clknet_leaf_139_clk_regs sg13g2_dfrbpq_1
X_05579_ net1197 net1212 _00000_ VPWR VGND sg13g2_nor2_1
X_07318_ net1246 net3759 net1150 _01029_ VPWR VGND sg13g2_mux2_1
X_08298_ net380 VGND VPWR net2096 i_exotiny._0031_\[0\] clknet_leaf_83_clk_regs sg13g2_dfrbpq_2
XFILLER_20_872 VPWR VGND sg13g2_fill_1
X_07249_ net2311 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[12\]
+ net1004 _00972_ VPWR VGND sg13g2_mux2_1
XFILLER_106_944 VPWR VGND sg13g2_decap_8
XFILLER_105_410 VPWR VGND sg13g2_decap_8
XFILLER_105_487 VPWR VGND sg13g2_decap_8
XFILLER_19_427 VPWR VGND sg13g2_fill_1
XFILLER_36_62 VPWR VGND sg13g2_fill_2
XFILLER_36_84 VPWR VGND sg13g2_decap_8
XFILLER_70_772 VPWR VGND sg13g2_fill_2
Xinput15 uio_in[5] net15 VPWR VGND sg13g2_buf_1
XFILLER_7_865 VPWR VGND sg13g2_fill_2
X_04950_ _01682_ _01680_ net1247 _01679_ _01421_ VPWR VGND sg13g2_a22oi_1
XFILLER_65_533 VPWR VGND sg13g2_fill_2
XFILLER_92_330 VPWR VGND sg13g2_decap_4
X_04881_ _01613_ net1258 VPWR VGND net1260 sg13g2_nand2b_2
X_06620_ net3155 net1155 _02670_ VPWR VGND sg13g2_nor2_1
X_08899__1083 VPWR VGND net1503 sg13g2_tiehi
X_06551_ VGND VPWR _01406_ net1216 _00620_ _02627_ sg13g2_a21oi_1
X_06482_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[13\]
+ net3019 net1025 _00563_ VPWR VGND sg13g2_mux2_1
X_05502_ _02194_ VPWR i_exotiny._1611_\[14\] VGND net1074 _02196_ sg13g2_o21ai_1
X_09270_ net81 VGND VPWR net2472 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[28\]
+ clknet_leaf_127_clk_regs sg13g2_dfrbpq_1
XFILLER_60_282 VPWR VGND sg13g2_fill_2
X_05433_ _02142_ _02128_ _02132_ VPWR VGND sg13g2_xnor2_1
X_08221_ net456 VGND VPWR _00302_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[20\]
+ clknet_leaf_172_clk_regs sg13g2_dfrbpq_1
XFILLER_20_102 VPWR VGND sg13g2_fill_2
X_05364_ _02086_ i_exotiny._2034_\[7\] _00021_ i_exotiny._2034_\[2\] _00016_ VPWR
+ VGND sg13g2_a22oi_1
X_08280__398 VPWR VGND net398 sg13g2_tiehi
X_08152_ net526 VGND VPWR net2221 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[16\]
+ clknet_leaf_131_clk_regs sg13g2_dfrbpq_1
X_08083_ net611 VGND VPWR net2235 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[20\]
+ clknet_leaf_86_clk_regs sg13g2_dfrbpq_1
X_07103_ net2936 _02943_ net913 _00856_ VPWR VGND sg13g2_mux2_1
X_05295_ _02021_ _01647_ i_exotiny._0032_\[0\] _01645_ i_exotiny._0025_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_07034_ net2410 i_exotiny._0017_\[0\] net1013 _00795_ VPWR VGND sg13g2_mux2_1
XFILLER_103_958 VPWR VGND sg13g2_decap_8
XFILLER_102_413 VPWR VGND sg13g2_decap_8
X_08686__1302 VPWR VGND net1722 sg13g2_tiehi
X_08985_ net1417 VGND VPWR net2027 i_exotiny._1160_\[6\] clknet_leaf_165_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_69_861 VPWR VGND sg13g2_fill_2
X_07936_ net712 VGND VPWR net1900 i_exotiny._1924_\[29\] clknet_leaf_30_clk_regs sg13g2_dfrbpq_1
XFILLER_57_28 VPWR VGND sg13g2_fill_2
XFILLER_69_883 VPWR VGND sg13g2_fill_1
XFILLER_68_360 VPWR VGND sg13g2_fill_2
X_07867_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[5\]
+ net2365 net978 _01334_ VPWR VGND sg13g2_mux2_1
X_08389__289 VPWR VGND net289 sg13g2_tiehi
X_06818_ VGND VPWR net3680 net1133 _02836_ _02835_ sg13g2_a21oi_1
X_07798_ net2935 net2869 net893 _01277_ VPWR VGND sg13g2_mux2_1
X_06749_ net3808 net1100 _02778_ VPWR VGND sg13g2_nor2_1
XFILLER_43_249 VPWR VGND sg13g2_fill_1
X_08506__174 VPWR VGND net174 sg13g2_tiehi
XFILLER_24_485 VPWR VGND sg13g2_fill_2
XFILLER_106_1028 VPWR VGND sg13g2_fill_1
X_08419_ net266 VGND VPWR _00493_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[18\]
+ clknet_leaf_90_clk_regs sg13g2_dfrbpq_1
XFILLER_22_75 VPWR VGND sg13g2_fill_1
XFILLER_4_813 VPWR VGND sg13g2_decap_8
XFILLER_3_312 VPWR VGND sg13g2_fill_2
XFILLER_106_741 VPWR VGND sg13g2_decap_8
XFILLER_3_334 VPWR VGND sg13g2_fill_1
XFILLER_105_284 VPWR VGND sg13g2_decap_8
Xfanout1113 _02091_ net1113 VPWR VGND sg13g2_buf_1
Xfanout1102 _02717_ net1102 VPWR VGND sg13g2_buf_8
Xfanout1124 net1125 net1124 VPWR VGND sg13g2_buf_8
Xfanout1135 net1136 net1135 VPWR VGND sg13g2_buf_8
X_08513__167 VPWR VGND net167 sg13g2_tiehi
Xfanout1146 _01484_ net1146 VPWR VGND sg13g2_buf_8
Xfanout1179 i_exotiny._0000_ net1179 VPWR VGND sg13g2_buf_8
Xfanout1157 net1158 net1157 VPWR VGND sg13g2_buf_8
Xfanout1168 _02414_ net1168 VPWR VGND sg13g2_buf_8
XFILLER_75_875 VPWR VGND sg13g2_fill_1
XFILLER_34_238 VPWR VGND sg13g2_fill_2
XFILLER_34_249 VPWR VGND sg13g2_fill_1
XFILLER_16_964 VPWR VGND sg13g2_fill_2
X_08764__1224 VPWR VGND net1644 sg13g2_tiehi
XFILLER_8_66 VPWR VGND sg13g2_fill_2
Xhold607 _00131_ VPWR VGND net2434 sg13g2_dlygate4sd3_1
Xhold618 _00141_ VPWR VGND net2445 sg13g2_dlygate4sd3_1
Xhold629 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[23\]
+ VPWR VGND net2456 sg13g2_dlygate4sd3_1
X_05080_ _01806_ _01811_ _01802_ _01812_ VPWR VGND sg13g2_nand3_1
XFILLER_98_923 VPWR VGND sg13g2_decap_8
XFILLER_97_422 VPWR VGND sg13g2_decap_8
Xhold2008 i_exotiny.i_wdg_top.o_wb_dat\[10\] VPWR VGND net3835 sg13g2_dlygate4sd3_1
X_07999__696 VPWR VGND net696 sg13g2_tiehi
XFILLER_100_917 VPWR VGND sg13g2_decap_8
Xhold1307 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[24\]
+ VPWR VGND net3134 sg13g2_dlygate4sd3_1
X_08095__599 VPWR VGND net599 sg13g2_tiehi
X_05982_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[8\]
+ net2154 net1050 _00184_ VPWR VGND sg13g2_mux2_1
Xhold1318 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[31\]
+ VPWR VGND net3145 sg13g2_dlygate4sd3_1
Xhold1329 _00647_ VPWR VGND net3156 sg13g2_dlygate4sd3_1
X_08770_ net1638 VGND VPWR net3369 i_exotiny._0015_\[1\] clknet_leaf_151_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_84_149 VPWR VGND sg13g2_fill_1
X_07721_ net2642 net2422 net995 _01217_ VPWR VGND sg13g2_mux2_1
X_04933_ _01665_ _01663_ _01664_ VPWR VGND sg13g2_nand2_1
XFILLER_65_352 VPWR VGND sg13g2_fill_2
X_07652_ net2396 net2888 net898 _01160_ VPWR VGND sg13g2_mux2_1
X_04864_ _01597_ net1266 _01446_ VPWR VGND sg13g2_nand2_1
X_07583_ _03159_ net3628 _01119_ VPWR VGND sg13g2_nor2_1
X_06603_ net1198 _02657_ _02658_ _00641_ VPWR VGND sg13g2_nor3_1
X_04795_ net1230 net1232 net1283 _01544_ VPWR VGND net3520 sg13g2_nand4_1
X_06534_ net2943 net2782 net930 _00609_ VPWR VGND sg13g2_mux2_1
X_09253_ net554 VGND VPWR _01308_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[11\]
+ clknet_leaf_130_clk_regs sg13g2_dfrbpq_1
X_06465_ net3064 net881 _02608_ _02611_ VPWR VGND sg13g2_mux2_1
X_09184_ net797 VGND VPWR _01239_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[6\]
+ clknet_leaf_79_clk_regs sg13g2_dfrbpq_1
X_05416_ VPWR i_exotiny._2043_\[9\] _02125_ VGND sg13g2_inv_1
X_08204_ net473 VGND VPWR net2116 i_exotiny._0037_\[3\] clknet_leaf_153_clk_regs sg13g2_dfrbpq_2
X_06396_ _02582_ _02581_ _01525_ _02180_ net3828 VPWR VGND sg13g2_a22oi_1
X_08135_ net1178 VGND VPWR net2013 _00023_ clknet_leaf_35_clk_regs sg13g2_dfrbpq_2
X_05347_ _02070_ net1116 _01578_ VPWR VGND sg13g2_nand2b_1
XFILLER_21_499 VPWR VGND sg13g2_fill_2
X_08066_ net628 VGND VPWR net3082 i_exotiny._0020_\[3\] clknet_leaf_84_clk_regs sg13g2_dfrbpq_2
X_05278_ VPWR VGND i_exotiny._0039_\[0\] _02003_ _01788_ i_exotiny._0033_\[0\] _02004_
+ _01772_ sg13g2_a221oi_1
Xclkbuf_leaf_118_clk_regs clknet_5_19__leaf_clk_regs clknet_leaf_118_clk_regs VPWR
+ VGND sg13g2_buf_8
X_07017_ net2746 net2994 net921 _00784_ VPWR VGND sg13g2_mux2_1
XFILLER_102_210 VPWR VGND sg13g2_decap_8
XFILLER_89_967 VPWR VGND sg13g2_decap_8
X_07939__709 VPWR VGND net709 sg13g2_tiehi
XFILLER_1_838 VPWR VGND sg13g2_decap_8
XFILLER_103_755 VPWR VGND sg13g2_decap_8
XFILLER_102_287 VPWR VGND sg13g2_decap_8
X_08968_ net1434 VGND VPWR net3769 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[4\]
+ clknet_leaf_14_clk_regs sg13g2_dfrbpq_1
XFILLER_84_650 VPWR VGND sg13g2_fill_2
X_07919_ net729 VGND VPWR net1923 i_exotiny._1924_\[12\] clknet_leaf_35_clk_regs sg13g2_dfrbpq_1
Xhold1841 i_exotiny._1619_\[0\] VPWR VGND net3668 sg13g2_dlygate4sd3_1
X_08899_ net1503 VGND VPWR _00957_ i_exotiny.i_wb_spi.dat_rx_r\[29\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_1
Xhold1852 i_exotiny._1489_\[1\] VPWR VGND net3679 sg13g2_dlygate4sd3_1
Xhold1863 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[3\] VPWR
+ VGND net3690 sg13g2_dlygate4sd3_1
Xhold1830 i_exotiny._6090_\[3\] VPWR VGND net3657 sg13g2_dlygate4sd3_1
Xhold1896 _03177_ VPWR VGND net3723 sg13g2_dlygate4sd3_1
Xhold1874 _01114_ VPWR VGND net3701 sg13g2_dlygate4sd3_1
XFILLER_17_706 VPWR VGND sg13g2_fill_2
X_08563__78 VPWR VGND net78 sg13g2_tiehi
XFILLER_29_566 VPWR VGND sg13g2_fill_1
Xhold1885 i_exotiny._1160_\[0\] VPWR VGND net3712 sg13g2_dlygate4sd3_1
XFILLER_17_42 VPWR VGND sg13g2_fill_1
XFILLER_44_525 VPWR VGND sg13g2_fill_1
XFILLER_24_293 VPWR VGND sg13g2_fill_1
X_08259__418 VPWR VGND net418 sg13g2_tiehi
XFILLER_4_698 VPWR VGND sg13g2_fill_2
XFILLER_95_926 VPWR VGND sg13g2_decap_8
Xhold4 _01115_ VPWR VGND net1831 sg13g2_dlygate4sd3_1
XFILLER_66_105 VPWR VGND sg13g2_fill_2
XFILLER_0_882 VPWR VGND sg13g2_decap_8
XFILLER_48_875 VPWR VGND sg13g2_fill_2
X_08818__1170 VPWR VGND net1590 sg13g2_tiehi
XFILLER_35_536 VPWR VGND sg13g2_decap_4
X_08166__512 VPWR VGND net512 sg13g2_tiehi
XFILLER_31_720 VPWR VGND sg13g2_fill_2
X_06250_ net2200 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[20\]
+ net1041 _00399_ VPWR VGND sg13g2_mux2_1
XFILLER_90_91 VPWR VGND sg13g2_fill_1
X_05201_ _01929_ _01780_ i_exotiny._0041_\[1\] _01761_ i_exotiny._0015_\[1\] VPWR
+ VGND sg13g2_a22oi_1
X_06181_ net2768 _02535_ net954 _00342_ VPWR VGND sg13g2_mux2_1
XFILLER_8_993 VPWR VGND sg13g2_decap_8
X_09282__57 VPWR VGND net57 sg13g2_tiehi
Xhold415 _01246_ VPWR VGND net2242 sg13g2_dlygate4sd3_1
Xhold404 _00348_ VPWR VGND net2231 sg13g2_dlygate4sd3_1
Xhold426 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[28\]
+ VPWR VGND net2253 sg13g2_dlygate4sd3_1
X_08379__299 VPWR VGND net299 sg13g2_tiehi
X_05132_ _01862_ _01780_ i_exotiny._0041_\[2\] _01778_ i_exotiny._0035_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold437 _00329_ VPWR VGND net2264 sg13g2_dlygate4sd3_1
Xhold448 _00589_ VPWR VGND net2275 sg13g2_dlygate4sd3_1
Xhold459 _00587_ VPWR VGND net2286 sg13g2_dlygate4sd3_1
X_05063_ _01795_ _01784_ i_exotiny._0042_\[3\] _01770_ i_exotiny._0025_\[3\] VPWR
+ VGND sg13g2_a22oi_1
Xfanout906 net907 net906 VPWR VGND sg13g2_buf_8
XFILLER_97_230 VPWR VGND sg13g2_fill_2
Xfanout939 net941 net939 VPWR VGND sg13g2_buf_8
Xfanout928 _02917_ net928 VPWR VGND sg13g2_buf_8
Xfanout917 _02941_ net917 VPWR VGND sg13g2_buf_8
X_08822_ net1586 VGND VPWR _00880_ i_exotiny.i_wb_spi.state_r\[21\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
Xhold1104 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[12\]
+ VPWR VGND net2931 sg13g2_dlygate4sd3_1
Xhold1115 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[19\]
+ VPWR VGND net2942 sg13g2_dlygate4sd3_1
X_08753_ net1655 VGND VPWR _00811_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[16\]
+ clknet_leaf_81_clk_regs sg13g2_dfrbpq_1
Xhold1137 i_exotiny._0026_\[3\] VPWR VGND net2964 sg13g2_dlygate4sd3_1
XFILLER_97_296 VPWR VGND sg13g2_decap_8
Xhold1148 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[19\]
+ VPWR VGND net2975 sg13g2_dlygate4sd3_1
X_05965_ i_exotiny._0020_\[1\] net884 _02486_ _02489_ VPWR VGND sg13g2_mux2_1
Xhold1126 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[17\]
+ VPWR VGND net2953 sg13g2_dlygate4sd3_1
Xhold1159 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[8\]
+ VPWR VGND net2986 sg13g2_dlygate4sd3_1
X_04916_ net1222 _01620_ _01640_ _01648_ VPWR VGND sg13g2_nor3_2
X_07704_ net2959 net3075 net996 _01200_ VPWR VGND sg13g2_mux2_1
X_05896_ i_exotiny._0019_\[1\] net2128 net977 _00113_ VPWR VGND sg13g2_mux2_1
XFILLER_65_182 VPWR VGND sg13g2_fill_1
X_08684_ net1724 VGND VPWR net3289 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[11\]
+ clknet_leaf_105_clk_regs sg13g2_dfrbpq_1
X_04847_ net1111 _01583_ _01585_ i_exotiny._1902_\[1\] VPWR VGND sg13g2_nor3_1
XFILLER_53_366 VPWR VGND sg13g2_decap_8
X_07635_ net2097 net2958 net899 _01143_ VPWR VGND sg13g2_mux2_1
X_07566_ _03147_ _03148_ _03149_ _01113_ VPWR VGND sg13g2_nor3_1
X_04778_ net1226 _01528_ _00012_ VPWR VGND sg13g2_nor2_1
X_06517_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[6\]
+ net2824 net929 _00592_ VPWR VGND sg13g2_mux2_1
X_09305_ net1353 VGND VPWR _01360_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[31\]
+ clknet_leaf_178_clk_regs sg13g2_dfrbpq_1
XFILLER_21_230 VPWR VGND sg13g2_fill_1
X_07497_ net3547 net3537 net905 _01080_ VPWR VGND sg13g2_mux2_1
X_09236_ net704 VGND VPWR _01291_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[26\]
+ clknet_leaf_135_clk_regs sg13g2_dfrbpq_1
X_08503__177 VPWR VGND net177 sg13g2_tiehi
X_06448_ net2381 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[13\]
+ net934 _00535_ VPWR VGND sg13g2_mux2_1
X_06379_ i_exotiny._0035_\[3\] net875 _02565_ _02570_ VPWR VGND sg13g2_mux2_1
X_09167_ net815 VGND VPWR net2388 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[23\]
+ clknet_leaf_173_clk_regs sg13g2_dfrbpq_1
X_09098_ net1304 VGND VPWR net2131 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[18\]
+ clknet_leaf_144_clk_regs sg13g2_dfrbpq_1
X_08118_ net576 VGND VPWR net2338 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[23\]
+ clknet_leaf_126_clk_regs sg13g2_dfrbpq_1
X_08049_ net645 VGND VPWR net2124 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[18\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
Xhold971 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[24\]
+ VPWR VGND net2798 sg13g2_dlygate4sd3_1
Xhold960 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[10\]
+ VPWR VGND net2787 sg13g2_dlygate4sd3_1
Xhold982 _01309_ VPWR VGND net2809 sg13g2_dlygate4sd3_1
Xhold993 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[23\]
+ VPWR VGND net2820 sg13g2_dlygate4sd3_1
XFILLER_88_263 VPWR VGND sg13g2_fill_1
XFILLER_0_189 VPWR VGND sg13g2_fill_1
Xhold1660 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[21\]
+ VPWR VGND net3487 sg13g2_dlygate4sd3_1
Xhold1671 i_exotiny._0314_\[15\] VPWR VGND net3498 sg13g2_dlygate4sd3_1
XFILLER_29_352 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_86_clk_regs clknet_5_31__leaf_clk_regs clknet_leaf_86_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_85_992 VPWR VGND sg13g2_decap_8
XFILLER_56_171 VPWR VGND sg13g2_fill_2
Xhold1693 i_exotiny._1715_ VPWR VGND net3520 sg13g2_dlygate4sd3_1
Xhold1682 i_exotiny._0314_\[12\] VPWR VGND net3509 sg13g2_dlygate4sd3_1
XFILLER_56_193 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_15_clk_regs clknet_5_6__leaf_clk_regs clknet_leaf_15_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_5_952 VPWR VGND sg13g2_decap_8
XFILLER_67_436 VPWR VGND sg13g2_fill_2
XFILLER_94_277 VPWR VGND sg13g2_decap_8
X_05750_ _02384_ net3634 _02383_ _00062_ VPWR VGND sg13g2_a21o_1
XFILLER_91_973 VPWR VGND sg13g2_decap_8
X_05681_ VGND VPWR i_exotiny._1616_\[0\] net1121 _02332_ _02331_ sg13g2_a21oi_1
X_04701_ net1224 _01458_ _01459_ VPWR VGND sg13g2_and2_1
X_07420_ i_exotiny._1160_\[17\] net1215 _03067_ VPWR VGND sg13g2_nor2_1
X_04632_ _01394_ net1257 VPWR VGND sg13g2_inv_2
XFILLER_50_347 VPWR VGND sg13g2_fill_2
X_07351_ net3307 _03009_ _03013_ VPWR VGND sg13g2_nor2b_1
X_06302_ net2814 net875 _02552_ _02557_ VPWR VGND sg13g2_mux2_1
X_07929__719 VPWR VGND net719 sg13g2_tiehi
XFILLER_31_561 VPWR VGND sg13g2_fill_2
X_07282_ net2202 net2789 net911 _00999_ VPWR VGND sg13g2_mux2_1
X_06233_ net2136 i_exotiny._0031_\[3\] net1039 _00382_ VPWR VGND sg13g2_mux2_1
X_09021_ net1381 VGND VPWR _01079_ i_exotiny._0315_\[9\] clknet_leaf_180_clk_regs
+ sg13g2_dfrbpq_1
Xhold201 i_exotiny.i_wdg_top.clk_div_inst.cnt\[7\] VPWR VGND net2028 sg13g2_dlygate4sd3_1
X_06164_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[12\]
+ net3245 net954 _00326_ VPWR VGND sg13g2_mux2_1
Xhold223 i_exotiny._1924_\[5\] VPWR VGND net2050 sg13g2_dlygate4sd3_1
X_08841__1145 VPWR VGND net1565 sg13g2_tiehi
Xhold212 _00648_ VPWR VGND net2039 sg13g2_dlygate4sd3_1
Xhold234 i_exotiny._0369_\[23\] VPWR VGND net2061 sg13g2_dlygate4sd3_1
X_05115_ _01844_ VPWR _01845_ VGND _01839_ _01843_ sg13g2_o21ai_1
XFILLER_105_839 VPWR VGND sg13g2_decap_8
XFILLER_104_327 VPWR VGND sg13g2_decap_8
Xhold278 i_exotiny.i_wb_spi.dat_rx_r\[10\] VPWR VGND net2105 sg13g2_dlygate4sd3_1
X_06095_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[21\]
+ net2593 net955 _00271_ VPWR VGND sg13g2_mux2_1
Xhold245 _01269_ VPWR VGND net2072 sg13g2_dlygate4sd3_1
Xhold256 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[28\]
+ VPWR VGND net2083 sg13g2_dlygate4sd3_1
Xhold267 _00766_ VPWR VGND net2094 sg13g2_dlygate4sd3_1
Xhold289 _00285_ VPWR VGND net2116 sg13g2_dlygate4sd3_1
X_05046_ net1220 _01754_ _01756_ _01778_ VPWR VGND sg13g2_nor3_2
XFILLER_100_500 VPWR VGND sg13g2_decap_8
X_08805_ net1603 VGND VPWR _00863_ i_exotiny.i_wb_spi.state_r\[4\] clknet_leaf_43_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_74_929 VPWR VGND sg13g2_fill_2
X_06997_ net3202 net3497 net920 _00764_ VPWR VGND sg13g2_mux2_1
XFILLER_85_299 VPWR VGND sg13g2_fill_1
X_05948_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[13\]
+ net2170 net969 _00157_ VPWR VGND sg13g2_mux2_1
X_08736_ net1672 VGND VPWR _00794_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[31\]
+ clknet_leaf_117_clk_regs sg13g2_dfrbpq_1
X_08249__428 VPWR VGND net428 sg13g2_tiehi
X_08667_ i_exotiny.i_wdg_top.cntr_inst.rst_n_sync VGND VPWR i_exotiny._2043_\[4\]
+ i_exotiny._2034_\[4\] net1229 sg13g2_dfrbpq_2
X_05879_ net5 _01473_ _02465_ VPWR VGND sg13g2_nor2_2
XFILLER_92_1019 VPWR VGND sg13g2_decap_8
X_07618_ net1205 net2055 _03182_ _01132_ VPWR VGND sg13g2_nor3_1
X_08598_ net1798 VGND VPWR _00670_ i_exotiny._1612_\[2\] clknet_leaf_28_clk_regs sg13g2_dfrbpq_2
XFILLER_26_399 VPWR VGND sg13g2_fill_2
XFILLER_42_859 VPWR VGND sg13g2_fill_1
X_07549_ net3658 _03137_ _03138_ VPWR VGND sg13g2_nor2_1
XFILLER_14_98 VPWR VGND sg13g2_fill_1
X_08792__1196 VPWR VGND net1616 sg13g2_tiehi
X_09219_ net760 VGND VPWR net2834 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[9\]
+ clknet_leaf_129_clk_regs sg13g2_dfrbpq_1
XFILLER_5_215 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_133_clk_regs clknet_5_20__leaf_clk_regs clknet_leaf_133_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08981__1001 VPWR VGND net1421 sg13g2_tiehi
XFILLER_100_2 VPWR VGND sg13g2_fill_1
XFILLER_2_922 VPWR VGND sg13g2_decap_8
Xhold790 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[28\]
+ VPWR VGND net2617 sg13g2_dlygate4sd3_1
X_08156__522 VPWR VGND net522 sg13g2_tiehi
XFILLER_103_360 VPWR VGND sg13g2_decap_8
XFILLER_49_414 VPWR VGND sg13g2_fill_2
XFILLER_2_999 VPWR VGND sg13g2_decap_8
XFILLER_36_108 VPWR VGND sg13g2_fill_1
XFILLER_45_620 VPWR VGND sg13g2_fill_2
Xhold1490 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[22\]
+ VPWR VGND net3317 sg13g2_dlygate4sd3_1
XFILLER_55_50 VPWR VGND sg13g2_fill_1
XFILLER_60_612 VPWR VGND sg13g2_fill_2
XFILLER_44_163 VPWR VGND sg13g2_fill_1
X_08163__515 VPWR VGND net515 sg13g2_tiehi
XFILLER_99_325 VPWR VGND sg13g2_decap_8
X_06920_ i_exotiny._0029_\[0\] net2635 net926 _00699_ VPWR VGND sg13g2_mux2_1
XFILLER_67_244 VPWR VGND sg13g2_fill_1
X_06851_ i_exotiny._0369_\[25\] net1189 _02863_ VPWR VGND sg13g2_nor2_1
XFILLER_83_759 VPWR VGND sg13g2_fill_2
XFILLER_83_726 VPWR VGND sg13g2_fill_1
X_06782_ VGND VPWR net1096 _02804_ _00673_ _02805_ sg13g2_a21oi_1
X_05802_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[1\] _02418_ net1262
+ _02419_ VPWR VGND sg13g2_nand3_1
X_05733_ _02370_ i_exotiny.i_wb_regs.spi_size_o\[0\] net1118 _02371_ VPWR VGND sg13g2_mux2_1
X_08521_ net159 VGND VPWR _00595_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[9\]
+ clknet_leaf_177_clk_regs sg13g2_dfrbpq_1
XFILLER_36_642 VPWR VGND sg13g2_decap_4
X_08452_ net228 VGND VPWR _00526_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[4\]
+ clknet_leaf_160_clk_regs sg13g2_dfrbpq_1
X_05664_ VGND VPWR i_exotiny._1617_\[0\] net1123 _02319_ _02318_ sg13g2_a21oi_1
XFILLER_51_656 VPWR VGND sg13g2_decap_8
X_08859__1127 VPWR VGND net1547 sg13g2_tiehi
XFILLER_23_347 VPWR VGND sg13g2_fill_1
XFILLER_24_848 VPWR VGND sg13g2_fill_2
X_07403_ net1079 net2022 _03054_ _01045_ VPWR VGND sg13g2_a21o_1
X_04615_ VPWR _01377_ net3511 VGND sg13g2_inv_1
XFILLER_51_678 VPWR VGND sg13g2_fill_1
X_08383_ net295 VGND VPWR _00464_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[21\]
+ clknet_leaf_139_clk_regs sg13g2_dfrbpq_1
X_05595_ _02267_ _01911_ _01909_ _02269_ VPWR VGND sg13g2_a21o_1
X_07334_ _02998_ _01404_ i_exotiny._0369_\[2\] VPWR VGND sg13g2_nand2_2
X_07265_ i_exotiny._0040_\[0\] net890 _02972_ _02974_ VPWR VGND sg13g2_mux2_1
X_06216_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[28\]
+ net2479 net948 _00371_ VPWR VGND sg13g2_mux2_1
X_09004_ net1398 VGND VPWR net3361 i_exotiny._1160_\[25\] clknet_leaf_162_clk_regs
+ sg13g2_dfrbpq_1
X_07196_ net3556 i_exotiny.i_wb_spi.dat_rx_r\[4\] net1093 _00932_ VPWR VGND sg13g2_mux2_1
XFILLER_105_636 VPWR VGND sg13g2_decap_8
X_06147_ net3442 net873 _02526_ _02531_ VPWR VGND sg13g2_mux2_1
XFILLER_104_124 VPWR VGND sg13g2_decap_8
X_06078_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[4\]
+ net3349 net957 _00254_ VPWR VGND sg13g2_mux2_1
X_08777__1211 VPWR VGND net1631 sg13g2_tiehi
XFILLER_99_870 VPWR VGND sg13g2_decap_8
X_05029_ net1238 net1240 net1237 _01761_ VGND VPWR _01754_ sg13g2_nor4_2
XFILLER_58_233 VPWR VGND sg13g2_fill_2
XFILLER_101_864 VPWR VGND sg13g2_decap_8
XFILLER_74_715 VPWR VGND sg13g2_fill_1
XFILLER_100_374 VPWR VGND sg13g2_decap_8
XFILLER_74_759 VPWR VGND sg13g2_fill_2
X_08700__1288 VPWR VGND net1708 sg13g2_tiehi
X_08719_ net1689 VGND VPWR _00777_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[14\]
+ clknet_leaf_123_clk_regs sg13g2_dfrbpq_1
XFILLER_42_634 VPWR VGND sg13g2_fill_2
XFILLER_25_64 VPWR VGND sg13g2_fill_1
XFILLER_6_524 VPWR VGND sg13g2_fill_1
XFILLER_97_807 VPWR VGND sg13g2_fill_1
XFILLER_49_211 VPWR VGND sg13g2_fill_1
XFILLER_2_796 VPWR VGND sg13g2_decap_8
X_07919__729 VPWR VGND net729 sg13g2_tiehi
Xclkbuf_leaf_30_clk_regs clknet_5_8__leaf_clk_regs clknet_leaf_30_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_2_46 VPWR VGND sg13g2_decap_4
XFILLER_32_122 VPWR VGND sg13g2_fill_1
X_05380_ VGND VPWR _02092_ _02097_ _02102_ _02101_ sg13g2_a21oi_1
X_07050_ net3255 net2393 net1014 _00811_ VPWR VGND sg13g2_mux2_1
X_06001_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[27\]
+ net2630 net1049 _00203_ VPWR VGND sg13g2_mux2_1
X_08239__438 VPWR VGND net438 sg13g2_tiehi
XFILLER_82_1018 VPWR VGND sg13g2_decap_8
X_07952_ net1179 VGND VPWR net3782 i_exotiny.i_wdg_top.do_cnt clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_2
X_06903_ _02904_ net3241 net3466 VPWR VGND sg13g2_nand2_1
XFILLER_96_851 VPWR VGND sg13g2_decap_8
X_07883_ net2981 net2810 net978 _01350_ VPWR VGND sg13g2_mux2_1
X_06834_ net1170 VPWR _02849_ VGND i_exotiny.i_wb_spi.dat_rx_r\[22\] net1185 sg13g2_o21ai_1
XFILLER_55_247 VPWR VGND sg13g2_fill_1
X_06765_ VGND VPWR _02788_ _02790_ _02791_ net1135 sg13g2_a21oi_1
X_08504_ net176 VGND VPWR _00578_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[24\]
+ clknet_leaf_108_clk_regs sg13g2_dfrbpq_1
XFILLER_55_269 VPWR VGND sg13g2_fill_1
XFILLER_37_995 VPWR VGND sg13g2_fill_1
X_05716_ net1114 net1899 _02358_ VPWR VGND sg13g2_nor2b_1
X_06696_ _02732_ net3741 _02725_ VPWR VGND sg13g2_nand2_1
X_05647_ net1125 net1922 _02306_ VPWR VGND sg13g2_nor2b_1
X_08435_ net250 VGND VPWR net3765 i_exotiny._0369_\[16\] clknet_leaf_16_clk_regs sg13g2_dfrbpq_2
X_08366_ net312 VGND VPWR _00447_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[4\]
+ clknet_leaf_139_clk_regs sg13g2_dfrbpq_1
X_05578_ net1204 i_exotiny._0000_ VPWR VGND sg13g2_inv_4
X_07317_ VGND VPWR _01404_ net1151 _01028_ _02985_ sg13g2_a21oi_1
X_08297_ net381 VGND VPWR net3209 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[31\]
+ clknet_leaf_99_clk_regs sg13g2_dfrbpq_1
X_07248_ net3352 net3386 net1006 _00971_ VPWR VGND sg13g2_mux2_1
XFILLER_106_923 VPWR VGND sg13g2_decap_8
X_07179_ _02126_ _02596_ _02953_ VPWR VGND sg13g2_nor2_1
XFILLER_105_466 VPWR VGND sg13g2_decap_8
X_08153__525 VPWR VGND net525 sg13g2_tiehi
XFILLER_98_1014 VPWR VGND sg13g2_decap_8
XFILLER_47_715 VPWR VGND sg13g2_decap_4
XFILLER_100_182 VPWR VGND sg13g2_fill_2
XFILLER_43_921 VPWR VGND sg13g2_fill_2
Xinput16 uio_in[6] net16 VPWR VGND sg13g2_buf_2
X_08160__518 VPWR VGND net518 sg13g2_tiehi
XFILLER_93_810 VPWR VGND sg13g2_fill_2
XFILLER_37_214 VPWR VGND sg13g2_fill_2
X_08269__409 VPWR VGND net409 sg13g2_tiehi
X_04880_ _01612_ _01609_ _01611_ VPWR VGND sg13g2_nand2_2
XFILLER_19_962 VPWR VGND sg13g2_fill_1
X_06550_ net1262 net1215 _02627_ VPWR VGND sg13g2_nor2_1
X_06481_ net3022 net3297 net1023 _00562_ VPWR VGND sg13g2_mux2_1
X_05501_ VGND VPWR net3407 net1276 _02196_ _02195_ sg13g2_a21oi_1
XFILLER_60_272 VPWR VGND sg13g2_fill_1
X_05432_ _02141_ _02140_ i_exotiny._1618_\[0\] _02135_ i_exotiny._1614_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_08220_ net457 VGND VPWR _00301_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[19\]
+ clknet_leaf_150_clk_regs sg13g2_dfrbpq_1
X_05363_ _02085_ _01399_ _01376_ _01398_ _01377_ VPWR VGND sg13g2_a22oi_1
X_08151_ net527 VGND VPWR net3061 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[15\]
+ clknet_leaf_118_clk_regs sg13g2_dfrbpq_1
X_08082_ net612 VGND VPWR _00163_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[19\]
+ clknet_leaf_92_clk_regs sg13g2_dfrbpq_1
X_07102_ i_exotiny._0015_\[1\] net881 _02940_ _02943_ VPWR VGND sg13g2_mux2_1
X_05294_ _02020_ _01653_ i_exotiny._0038_\[0\] _01642_ i_exotiny._0015_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_07033_ VGND VPWR net1166 _02935_ _02934_ net1139 sg13g2_a21oi_2
XFILLER_103_937 VPWR VGND sg13g2_decap_8
X_08984_ net1418 VGND VPWR net1997 i_exotiny._1160_\[5\] clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
XFILLER_102_469 VPWR VGND sg13g2_decap_8
X_07935_ net713 VGND VPWR net1919 i_exotiny._1924_\[28\] clknet_leaf_30_clk_regs sg13g2_dfrbpq_1
X_08575__54 VPWR VGND net54 sg13g2_tiehi
X_07866_ net2069 net2684 net982 _01333_ VPWR VGND sg13g2_mux2_1
XFILLER_84_898 VPWR VGND sg13g2_fill_2
X_06817_ net1132 _02833_ _02834_ _02835_ VPWR VGND sg13g2_nor3_1
X_07797_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[11\]
+ net2251 net891 _01276_ VPWR VGND sg13g2_mux2_1
XFILLER_44_707 VPWR VGND sg13g2_fill_1
X_06748_ VGND VPWR net2042 net1130 _02777_ _02776_ sg13g2_a21oi_1
XFILLER_12_604 VPWR VGND sg13g2_fill_2
XFILLER_40_913 VPWR VGND sg13g2_fill_2
XFILLER_106_1007 VPWR VGND sg13g2_decap_8
X_08418_ net267 VGND VPWR _00492_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[17\]
+ clknet_leaf_90_clk_regs sg13g2_dfrbpq_1
X_06679_ _01362_ _02712_ _02716_ VPWR VGND sg13g2_nor2_1
X_08349_ net329 VGND VPWR net2821 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[19\]
+ clknet_leaf_98_clk_regs sg13g2_dfrbpq_1
X_07909__739 VPWR VGND net739 sg13g2_tiehi
XFILLER_106_720 VPWR VGND sg13g2_decap_8
XFILLER_4_869 VPWR VGND sg13g2_decap_8
XFILLER_106_797 VPWR VGND sg13g2_decap_8
XFILLER_105_263 VPWR VGND sg13g2_decap_8
Xfanout1103 net1104 net1103 VPWR VGND sg13g2_buf_2
Xfanout1125 _01582_ net1125 VPWR VGND sg13g2_buf_8
Xfanout1114 net1115 net1114 VPWR VGND sg13g2_buf_2
Xfanout1147 _03050_ net1147 VPWR VGND sg13g2_buf_8
Xfanout1136 _01507_ net1136 VPWR VGND sg13g2_buf_2
Xfanout1169 _01517_ net1169 VPWR VGND sg13g2_buf_8
X_08854__1132 VPWR VGND net1552 sg13g2_tiehi
Xfanout1158 _02415_ net1158 VPWR VGND sg13g2_buf_8
XFILLER_35_707 VPWR VGND sg13g2_fill_2
XFILLER_90_857 VPWR VGND sg13g2_fill_2
X_08229__448 VPWR VGND net448 sg13g2_tiehi
X_09279__63 VPWR VGND net63 sg13g2_tiehi
X_07982__123 VPWR VGND net123 sg13g2_tiehi
Xhold608 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[27\]
+ VPWR VGND net2435 sg13g2_dlygate4sd3_1
Xhold619 i_exotiny._0314_\[28\] VPWR VGND net2446 sg13g2_dlygate4sd3_1
XFILLER_98_902 VPWR VGND sg13g2_decap_8
XFILLER_97_401 VPWR VGND sg13g2_decap_8
XFILLER_40_4 VPWR VGND sg13g2_fill_1
Xhold2009 i_exotiny._0079_\[1\] VPWR VGND net3836 sg13g2_dlygate4sd3_1
XFILLER_98_979 VPWR VGND sg13g2_decap_8
XFILLER_97_467 VPWR VGND sg13g2_decap_4
XFILLER_2_390 VPWR VGND sg13g2_fill_1
Xhold1308 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[27\]
+ VPWR VGND net3135 sg13g2_dlygate4sd3_1
Xhold1319 _01166_ VPWR VGND net3146 sg13g2_dlygate4sd3_1
X_07720_ net2748 net3079 net994 _01216_ VPWR VGND sg13g2_mux2_1
X_08557__98 VPWR VGND net98 sg13g2_tiehi
XFILLER_38_501 VPWR VGND sg13g2_fill_1
X_05981_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[7\]
+ net2440 net1051 _00183_ VPWR VGND sg13g2_mux2_1
XFILLER_93_640 VPWR VGND sg13g2_fill_2
X_04932_ _01664_ _01630_ i_exotiny._0041_\[3\] _01626_ i_exotiny._0014_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_04863_ _01596_ VPWR i_exotiny._1902_\[6\] VGND _01580_ _01595_ sg13g2_o21ai_1
X_07651_ net2236 net3085 net899 _01159_ VPWR VGND sg13g2_mux2_1
XFILLER_38_589 VPWR VGND sg13g2_fill_2
X_07582_ net1179 VPWR _03160_ VGND net3627 _03158_ sg13g2_o21ai_1
X_08388__290 VPWR VGND net290 sg13g2_tiehi
X_06602_ net2864 net1154 _02658_ VPWR VGND sg13g2_nor2_1
X_09236__704 VPWR VGND net704 sg13g2_tiehi
X_04794_ _01543_ net1283 net3702 VPWR VGND sg13g2_nand2_1
X_06533_ net2437 net2965 net929 _00608_ VPWR VGND sg13g2_mux2_1
X_06464_ _02610_ net3328 net938 _00550_ VPWR VGND sg13g2_mux2_1
X_09252_ net555 VGND VPWR net2143 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[10\]
+ clknet_leaf_126_clk_regs sg13g2_dfrbpq_1
X_09183_ net798 VGND VPWR _01238_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[5\]
+ clknet_leaf_80_clk_regs sg13g2_dfrbpq_1
X_05415_ _02124_ VPWR _02125_ VGND i_exotiny._2034_\[9\] _02123_ sg13g2_o21ai_1
X_06395_ i_exotiny._0315_\[8\] net3476 net1272 _02581_ VPWR VGND sg13g2_mux2_1
X_08203_ net474 VGND VPWR net2962 i_exotiny._0037_\[2\] clknet_leaf_152_clk_regs sg13g2_dfrbpq_2
X_08397__537 VPWR VGND net537 sg13g2_tiehi
X_08134_ net1177 VGND VPWR net2064 _00022_ clknet_leaf_35_clk_regs sg13g2_dfrbpq_2
X_05346_ VGND VPWR i_exotiny._1207_ _02069_ _02055_ sg13g2_or2_1
X_08065_ net629 VGND VPWR net2169 i_exotiny._0020_\[2\] clknet_leaf_85_clk_regs sg13g2_dfrbpq_2
X_05277_ _01989_ _02001_ _01755_ _02003_ VPWR VGND _02002_ sg13g2_nand4_1
XFILLER_1_817 VPWR VGND sg13g2_decap_8
X_07016_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[20\]
+ net3395 net922 _00783_ VPWR VGND sg13g2_mux2_1
XFILLER_103_734 VPWR VGND sg13g2_decap_8
XFILLER_89_946 VPWR VGND sg13g2_decap_8
X_08635__1342 VPWR VGND net1762 sg13g2_tiehi
XFILLER_102_266 VPWR VGND sg13g2_decap_8
XFILLER_75_117 VPWR VGND sg13g2_fill_2
XFILLER_29_501 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_158_clk_regs clknet_5_18__leaf_clk_regs clknet_leaf_158_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08967_ net1435 VGND VPWR net3691 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[3\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
Xhold1820 i_exotiny._0369_\[24\] VPWR VGND net3647 sg13g2_dlygate4sd3_1
Xhold1831 i_exotiny.i_rstctl.cnt\[3\] VPWR VGND net3658 sg13g2_dlygate4sd3_1
X_07918_ net730 VGND VPWR net1910 i_exotiny._1924_\[11\] clknet_leaf_34_clk_regs sg13g2_dfrbpq_1
Xhold1853 i_exotiny._1617_\[3\] VPWR VGND net3680 sg13g2_dlygate4sd3_1
Xhold1842 _00688_ VPWR VGND net3669 sg13g2_dlygate4sd3_1
X_08898_ net1504 VGND VPWR _00956_ i_exotiny.i_wb_spi.dat_rx_r\[28\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_1
X_08150__528 VPWR VGND net528 sg13g2_tiehi
Xhold1886 i_exotiny.i_wb_qspi_mem.cnt_r\[2\] VPWR VGND net3713 sg13g2_dlygate4sd3_1
Xhold1875 i_exotiny._1711_ VPWR VGND net3702 sg13g2_dlygate4sd3_1
X_07849_ net2910 net3273 net983 _01322_ VPWR VGND sg13g2_mux2_1
Xhold1864 _01025_ VPWR VGND net3691 sg13g2_dlygate4sd3_1
XFILLER_95_1028 VPWR VGND sg13g2_fill_1
XFILLER_95_1017 VPWR VGND sg13g2_decap_8
Xhold1897 i_exotiny._1725_ VPWR VGND net3724 sg13g2_dlygate4sd3_1
XFILLER_71_356 VPWR VGND sg13g2_fill_2
X_08443__240 VPWR VGND net240 sg13g2_tiehi
XFILLER_13_913 VPWR VGND sg13g2_fill_1
XFILLER_9_939 VPWR VGND sg13g2_decap_8
XFILLER_106_594 VPWR VGND sg13g2_decap_8
XFILLER_95_905 VPWR VGND sg13g2_decap_8
XFILLER_0_861 VPWR VGND sg13g2_decap_8
Xhold5 i_exotiny.i_wdg_top.fsm_inst.sw_trg_s1wto VPWR VGND net1832 sg13g2_dlygate4sd3_1
XFILLER_59_180 VPWR VGND sg13g2_fill_1
XFILLER_47_342 VPWR VGND sg13g2_fill_1
XFILLER_62_312 VPWR VGND sg13g2_fill_2
XFILLER_15_283 VPWR VGND sg13g2_fill_2
Xclkbuf_4_2_0_clk_regs clknet_0_clk_regs clknet_4_2_0_clk_regs VPWR VGND sg13g2_buf_8
X_08713__1275 VPWR VGND net1695 sg13g2_tiehi
X_05200_ _01928_ _01787_ i_exotiny._0031_\[1\] _01776_ i_exotiny._0021_\[1\] VPWR
+ VGND sg13g2_a22oi_1
X_06180_ net890 net3269 _02533_ _02535_ VPWR VGND sg13g2_mux2_1
XFILLER_8_972 VPWR VGND sg13g2_decap_8
Xhold416 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[6\]
+ VPWR VGND net2243 sg13g2_dlygate4sd3_1
Xhold427 _01353_ VPWR VGND net2254 sg13g2_dlygate4sd3_1
Xhold405 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[9\]
+ VPWR VGND net2232 sg13g2_dlygate4sd3_1
X_05131_ VPWR VGND i_exotiny._0031_\[2\] _01860_ _01787_ i_exotiny._0020_\[2\] _01861_
+ _01779_ sg13g2_a221oi_1
XFILLER_104_509 VPWR VGND sg13g2_decap_8
Xhold449 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[28\]
+ VPWR VGND net2276 sg13g2_dlygate4sd3_1
Xhold438 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[17\]
+ VPWR VGND net2265 sg13g2_dlygate4sd3_1
X_05062_ _01794_ _01790_ i_exotiny._0034_\[3\] _01780_ i_exotiny._0041_\[3\] VPWR
+ VGND sg13g2_a22oi_1
Xfanout907 _03105_ net907 VPWR VGND sg13g2_buf_8
X_08821_ net1587 VGND VPWR _00879_ i_exotiny.i_wb_spi.state_r\[20\] clknet_leaf_41_clk_regs
+ sg13g2_dfrbpq_1
Xfanout929 net931 net929 VPWR VGND sg13g2_buf_8
XFILLER_31_0 VPWR VGND sg13g2_decap_8
Xfanout918 net923 net918 VPWR VGND sg13g2_buf_8
XFILLER_97_275 VPWR VGND sg13g2_decap_8
Xhold1105 _00120_ VPWR VGND net2932 sg13g2_dlygate4sd3_1
X_08935__1047 VPWR VGND net1467 sg13g2_tiehi
X_07938__710 VPWR VGND net710 sg13g2_tiehi
X_08752_ net1656 VGND VPWR net3200 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[15\]
+ clknet_leaf_87_clk_regs sg13g2_dfrbpq_1
Xhold1127 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[15\]
+ VPWR VGND net2954 sg13g2_dlygate4sd3_1
X_05964_ net2812 _02488_ net968 _00172_ VPWR VGND sg13g2_mux2_1
Xhold1116 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[23\]
+ VPWR VGND net2943 sg13g2_dlygate4sd3_1
Xhold1138 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[26\]
+ VPWR VGND net2965 sg13g2_dlygate4sd3_1
Xhold1149 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[28\]
+ VPWR VGND net2976 sg13g2_dlygate4sd3_1
X_08683_ net1725 VGND VPWR net3217 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[10\]
+ clknet_leaf_104_clk_regs sg13g2_dfrbpq_1
X_07703_ net2992 i_exotiny._0027_\[0\] net994 _01199_ VPWR VGND sg13g2_mux2_1
X_04915_ net1259 net1261 net1223 _01647_ VGND VPWR _01640_ sg13g2_nor4_2
X_05895_ i_exotiny._0019_\[0\] net2482 net975 _00112_ VPWR VGND sg13g2_mux2_1
X_07634_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[7\]
+ net2859 net896 _01142_ VPWR VGND sg13g2_mux2_1
X_04846_ net3728 net1840 _01585_ VPWR VGND sg13g2_xor2_1
X_04777_ _01525_ _01527_ _01528_ VPWR VGND sg13g2_nor2_1
X_07565_ _03149_ net1283 _01486_ VPWR VGND sg13g2_nand2_1
XFILLER_22_710 VPWR VGND sg13g2_fill_1
X_06516_ net2285 net2541 net932 _00591_ VPWR VGND sg13g2_mux2_1
X_09304_ net1355 VGND VPWR net3067 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[30\]
+ clknet_leaf_171_clk_regs sg13g2_dfrbpq_1
X_07496_ net3545 net3555 net904 _01079_ VPWR VGND sg13g2_mux2_1
X_06447_ net2737 net3003 net937 _00534_ VPWR VGND sg13g2_mux2_1
XFILLER_21_242 VPWR VGND sg13g2_fill_1
X_09235_ net744 VGND VPWR net2681 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[25\]
+ clknet_leaf_130_clk_regs sg13g2_dfrbpq_1
XFILLER_10_949 VPWR VGND sg13g2_decap_8
X_06378_ _02569_ net2718 net1030 _00505_ VPWR VGND sg13g2_mux2_1
X_09166_ net816 VGND VPWR _01221_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[22\]
+ clknet_leaf_172_clk_regs sg13g2_dfrbpq_1
X_08117_ net577 VGND VPWR net3265 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[22\]
+ clknet_leaf_122_clk_regs sg13g2_dfrbpq_1
X_09097_ net1305 VGND VPWR net3312 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[17\]
+ clknet_leaf_143_clk_regs sg13g2_dfrbpq_1
X_05329_ i_exotiny._0352_ _01817_ _02053_ VPWR VGND sg13g2_nor2_1
X_08048_ net646 VGND VPWR net2490 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[17\]
+ clknet_leaf_55_clk_regs sg13g2_dfrbpq_1
Xhold972 _00270_ VPWR VGND net2799 sg13g2_dlygate4sd3_1
Xhold950 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[6\]
+ VPWR VGND net2777 sg13g2_dlygate4sd3_1
Xhold961 _00901_ VPWR VGND net2788 sg13g2_dlygate4sd3_1
XFILLER_103_542 VPWR VGND sg13g2_decap_4
Xhold994 _00430_ VPWR VGND net2821 sg13g2_dlygate4sd3_1
Xhold983 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[25\]
+ VPWR VGND net2810 sg13g2_dlygate4sd3_1
X_08219__458 VPWR VGND net458 sg13g2_tiehi
XFILLER_95_48 VPWR VGND sg13g2_fill_2
Xhold1650 _00632_ VPWR VGND net3477 sg13g2_dlygate4sd3_1
Xhold1661 _00193_ VPWR VGND net3488 sg13g2_dlygate4sd3_1
Xhold1683 i_exotiny._0033_\[3\] VPWR VGND net3510 sg13g2_dlygate4sd3_1
XFILLER_56_150 VPWR VGND sg13g2_fill_1
Xhold1694 _01494_ VPWR VGND net3521 sg13g2_dlygate4sd3_1
Xhold1672 _00639_ VPWR VGND net3499 sg13g2_dlygate4sd3_1
XFILLER_44_323 VPWR VGND sg13g2_fill_2
XFILLER_72_654 VPWR VGND sg13g2_fill_2
XFILLER_44_52 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_55_clk_regs clknet_5_15__leaf_clk_regs clknet_leaf_55_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_12_297 VPWR VGND sg13g2_fill_1
XFILLER_60_62 VPWR VGND sg13g2_fill_1
XFILLER_8_268 VPWR VGND sg13g2_fill_2
XFILLER_5_931 VPWR VGND sg13g2_decap_8
XFILLER_99_507 VPWR VGND sg13g2_decap_8
XFILLER_106_391 VPWR VGND sg13g2_decap_8
XFILLER_54_109 VPWR VGND sg13g2_fill_1
X_04700_ net1251 net1252 _01456_ _01458_ VPWR VGND sg13g2_nor3_1
XFILLER_91_952 VPWR VGND sg13g2_decap_8
X_05680_ net1121 i_exotiny._1924_\[20\] _02331_ VPWR VGND sg13g2_nor2b_1
X_08385__293 VPWR VGND net293 sg13g2_tiehi
XFILLER_35_378 VPWR VGND sg13g2_fill_2
X_04631_ net3784 _01393_ VPWR VGND sg13g2_inv_4
X_07350_ net3727 net1078 _03012_ VPWR VGND sg13g2_nor2_1
X_06301_ _02556_ net3206 net939 _00441_ VPWR VGND sg13g2_mux2_1
X_07281_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[6\]
+ net2584 net909 _00998_ VPWR VGND sg13g2_mux2_1
X_09020_ net1382 VGND VPWR _01078_ i_exotiny._0315_\[8\] clknet_leaf_3_clk_regs sg13g2_dfrbpq_2
XFILLER_102_1021 VPWR VGND sg13g2_decap_8
X_06232_ net3336 net3231 net1041 _00381_ VPWR VGND sg13g2_mux2_1
Xhold202 _03164_ VPWR VGND net2029 sg13g2_dlygate4sd3_1
X_06163_ net2739 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[15\]
+ net950 _00325_ VPWR VGND sg13g2_mux2_1
XFILLER_105_818 VPWR VGND sg13g2_decap_8
XFILLER_85_1027 VPWR VGND sg13g2_fill_2
Xhold224 _00030_ VPWR VGND net2051 sg13g2_dlygate4sd3_1
Xhold235 i_exotiny._1611_\[19\] VPWR VGND net2062 sg13g2_dlygate4sd3_1
Xhold213 i_exotiny._1160_\[14\] VPWR VGND net2040 sg13g2_dlygate4sd3_1
X_05114_ VGND VPWR net1267 i_exotiny._6090_\[2\] _01844_ _01750_ sg13g2_a21oi_1
XFILLER_104_306 VPWR VGND sg13g2_decap_8
Xhold268 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[4\]
+ VPWR VGND net2095 sg13g2_dlygate4sd3_1
Xhold246 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[19\]
+ VPWR VGND net2073 sg13g2_dlygate4sd3_1
X_06094_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[20\]
+ net2798 net956 _00270_ VPWR VGND sg13g2_mux2_1
Xhold257 _00787_ VPWR VGND net2084 sg13g2_dlygate4sd3_1
Xhold279 i_exotiny.i_wb_regs.spi_cpol_o VPWR VGND net2106 sg13g2_dlygate4sd3_1
X_08392__286 VPWR VGND net286 sg13g2_tiehi
X_05045_ net1235 _01756_ _01759_ _01777_ VPWR VGND sg13g2_nor3_2
X_08804_ net1604 VGND VPWR _00862_ i_exotiny.i_wb_spi.state_r\[3\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_58_437 VPWR VGND sg13g2_fill_2
X_06996_ i_exotiny._0032_\[0\] net2059 net922 _00763_ VPWR VGND sg13g2_mux2_1
X_08735_ net1673 VGND VPWR net3078 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[30\]
+ clknet_leaf_116_clk_regs sg13g2_dfrbpq_1
X_05947_ net2792 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[16\]
+ net968 _00156_ VPWR VGND sg13g2_mux2_1
XFILLER_45_109 VPWR VGND sg13g2_fill_2
X_08666_ net1203 VGND VPWR i_exotiny._2043_\[3\] i_exotiny._2034_\[3\] net1228 sg13g2_dfrbpq_2
XFILLER_82_952 VPWR VGND sg13g2_fill_2
X_05878_ _02464_ net2891 net1055 _00110_ VPWR VGND sg13g2_mux2_1
XFILLER_54_665 VPWR VGND sg13g2_fill_2
X_04829_ _01567_ _01568_ _01566_ _01569_ VPWR VGND sg13g2_nand3_1
X_07617_ net2054 _03180_ _03182_ VPWR VGND sg13g2_and2_1
X_08597_ net1799 VGND VPWR _00669_ i_exotiny._1612_\[1\] clknet_leaf_31_clk_regs sg13g2_dfrbpq_2
X_08585__1392 VPWR VGND net1812 sg13g2_tiehi
X_07548_ _03133_ net2299 _03137_ _01107_ VPWR VGND sg13g2_nor3_1
XFILLER_41_348 VPWR VGND sg13g2_fill_1
X_07479_ VPWR _03106_ net902 VGND sg13g2_inv_1
X_09218_ net761 VGND VPWR _01273_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[8\]
+ clknet_leaf_136_clk_regs sg13g2_dfrbpq_1
X_09149_ net833 VGND VPWR _01204_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[5\]
+ clknet_leaf_172_clk_regs sg13g2_dfrbpq_1
X_08809__1179 VPWR VGND net1599 sg13g2_tiehi
XFILLER_1_400 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_173_clk_regs clknet_5_5__leaf_clk_regs clknet_leaf_173_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_2_901 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_102_clk_regs clknet_5_23__leaf_clk_regs clknet_leaf_102_clk_regs VPWR
+ VGND sg13g2_buf_8
Xhold791 _00610_ VPWR VGND net2618 sg13g2_dlygate4sd3_1
Xhold780 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[9\]
+ VPWR VGND net2607 sg13g2_dlygate4sd3_1
XFILLER_77_702 VPWR VGND sg13g2_fill_2
XFILLER_49_404 VPWR VGND sg13g2_fill_1
XFILLER_2_978 VPWR VGND sg13g2_decap_8
XFILLER_104_895 VPWR VGND sg13g2_decap_8
XFILLER_92_716 VPWR VGND sg13g2_fill_1
Xhold1491 i_exotiny._0315_\[21\] VPWR VGND net3318 sg13g2_dlygate4sd3_1
Xhold1480 i_exotiny._0369_\[22\] VPWR VGND net3307 sg13g2_dlygate4sd3_1
XFILLER_44_120 VPWR VGND sg13g2_decap_8
X_07928__720 VPWR VGND net720 sg13g2_tiehi
XFILLER_99_304 VPWR VGND sg13g2_decap_8
XFILLER_5_783 VPWR VGND sg13g2_decap_4
X_06850_ VGND VPWR net1094 _02861_ _00684_ _02862_ sg13g2_a21oi_1
X_07935__713 VPWR VGND net713 sg13g2_tiehi
X_05801_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[0\] _02417_ _02418_
+ VPWR VGND sg13g2_and2_1
X_06781_ net3559 net1096 _02805_ VPWR VGND sg13g2_nor2_1
XFILLER_64_930 VPWR VGND sg13g2_fill_2
XFILLER_48_470 VPWR VGND sg13g2_fill_2
X_05732_ _02370_ net1972 _02367_ VPWR VGND sg13g2_xnor2_1
X_09289__1401 VPWR VGND net1821 sg13g2_tiehi
X_08520_ net160 VGND VPWR net3154 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[8\]
+ clknet_leaf_176_clk_regs sg13g2_dfrbpq_1
X_05663_ net1122 net2004 _02318_ VPWR VGND sg13g2_nor2b_1
XFILLER_51_613 VPWR VGND sg13g2_fill_2
XFILLER_35_142 VPWR VGND sg13g2_fill_1
X_08451_ net229 VGND VPWR net3345 i_exotiny._0039_\[3\] clknet_leaf_157_clk_regs sg13g2_dfrbpq_2
X_04614_ VPWR _01376_ _00015_ VGND sg13g2_inv_1
XFILLER_51_635 VPWR VGND sg13g2_decap_8
X_07402_ net1079 _03049_ _03053_ _03054_ VPWR VGND sg13g2_nor3_1
X_08885__1097 VPWR VGND net1517 sg13g2_tiehi
X_08382_ net296 VGND VPWR _00463_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[20\]
+ clknet_leaf_138_clk_regs sg13g2_dfrbpq_1
X_05594_ VGND VPWR _01911_ _02267_ _02268_ _01909_ sg13g2_a21oi_1
X_08209__468 VPWR VGND net468 sg13g2_tiehi
X_07333_ _02997_ i_exotiny._0369_\[4\] i_exotiny._0369_\[5\] VPWR VGND sg13g2_nand2_1
X_07264_ net3173 net2542 net1006 _00987_ VPWR VGND sg13g2_mux2_1
X_06215_ net2717 net2475 net947 _00370_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_0_clk_regs clknet_5_0__leaf_clk_regs clknet_leaf_0_clk_regs VPWR VGND
+ sg13g2_buf_8
X_09003_ net1399 VGND VPWR net3385 i_exotiny._1160_\[24\] clknet_leaf_17_clk_regs
+ sg13g2_dfrbpq_1
X_07195_ net3574 net3556 net1093 _00931_ VPWR VGND sg13g2_mux2_1
XFILLER_3_709 VPWR VGND sg13g2_fill_1
XFILLER_105_615 VPWR VGND sg13g2_decap_8
X_06146_ _02530_ net2664 net1045 _00312_ VPWR VGND sg13g2_mux2_1
X_08255__422 VPWR VGND net422 sg13g2_tiehi
X_06077_ i_exotiny._0038_\[3\] net2303 net960 _00253_ VPWR VGND sg13g2_mux2_1
X_05028_ net1235 _01753_ _01759_ _01760_ VPWR VGND sg13g2_nor3_2
XFILLER_101_843 VPWR VGND sg13g2_decap_8
XFILLER_100_353 VPWR VGND sg13g2_decap_8
XFILLER_86_576 VPWR VGND sg13g2_fill_2
XFILLER_47_908 VPWR VGND sg13g2_fill_2
X_06979_ net1994 net2656 net1018 _00752_ VPWR VGND sg13g2_mux2_1
XFILLER_27_643 VPWR VGND sg13g2_fill_1
X_08718_ net1690 VGND VPWR net2076 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[13\]
+ clknet_leaf_120_clk_regs sg13g2_dfrbpq_1
XFILLER_82_782 VPWR VGND sg13g2_fill_2
X_08649_ net1748 VGND VPWR net2279 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[18\]
+ clknet_leaf_149_clk_regs sg13g2_dfrbpq_1
XFILLER_26_175 VPWR VGND sg13g2_fill_1
X_08262__415 VPWR VGND net415 sg13g2_tiehi
XFILLER_42_668 VPWR VGND sg13g2_fill_2
X_08930__1052 VPWR VGND net1472 sg13g2_tiehi
XFILLER_9_0 VPWR VGND sg13g2_fill_1
XFILLER_2_775 VPWR VGND sg13g2_decap_8
XFILLER_104_692 VPWR VGND sg13g2_decap_8
XFILLER_96_329 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_106_90 VPWR VGND sg13g2_decap_8
XFILLER_66_61 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_70_clk_regs clknet_5_25__leaf_clk_regs clknet_leaf_70_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_17_131 VPWR VGND sg13g2_fill_1
X_08382__296 VPWR VGND net296 sg13g2_tiehi
XFILLER_32_189 VPWR VGND sg13g2_fill_1
XFILLER_41_690 VPWR VGND sg13g2_decap_8
X_08278__400 VPWR VGND net400 sg13g2_tiehi
X_06000_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[26\]
+ net2156 net1048 _00202_ VPWR VGND sg13g2_mux2_1
X_08750__1238 VPWR VGND net1658 sg13g2_tiehi
X_07951_ net95 VGND VPWR net1932 i_exotiny.i_wb_spi.cnt_hbit_r\[6\] clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_1
X_06902_ net3658 net2298 net3681 _02902_ _02903_ VPWR VGND sg13g2_nor4_1
X_07882_ net2327 net2412 net979 _01349_ VPWR VGND sg13g2_mux2_1
X_06833_ net3307 net1188 _02848_ VPWR VGND sg13g2_nor2_1
X_06764_ _02789_ VPWR _02790_ VGND net3641 net1190 sg13g2_o21ai_1
X_09299__1119 VPWR VGND net1539 sg13g2_tiehi
X_08503_ net177 VGND VPWR _00577_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[23\]
+ clknet_leaf_109_clk_regs sg13g2_dfrbpq_1
X_05715_ net1998 net1059 _02357_ VPWR VGND sg13g2_nor2_1
XFILLER_52_955 VPWR VGND sg13g2_fill_2
XFILLER_51_421 VPWR VGND sg13g2_fill_2
X_06695_ VPWR VGND _01506_ _02731_ _02730_ _01361_ _00660_ _02719_ sg13g2_a221oi_1
X_05646_ VGND VPWR net1066 _02305_ _00037_ _02303_ sg13g2_a21oi_1
XFILLER_23_134 VPWR VGND sg13g2_fill_2
X_08434_ net251 VGND VPWR _00508_ i_exotiny._0369_\[28\] clknet_leaf_16_clk_regs sg13g2_dfrbpq_2
X_05577_ _02256_ net2570 net1291 VPWR VGND sg13g2_nand2_1
X_08365_ net313 VGND VPWR _00446_ i_exotiny._0014_\[3\] clknet_leaf_141_clk_regs sg13g2_dfrbpq_2
X_07316_ net3684 net1150 _02985_ VPWR VGND sg13g2_nor2_1
X_08296_ net382 VGND VPWR net2672 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[30\]
+ clknet_leaf_106_clk_regs sg13g2_dfrbpq_1
X_07247_ net2487 net2361 net1003 _00970_ VPWR VGND sg13g2_mux2_1
XFILLER_106_902 VPWR VGND sg13g2_decap_8
XFILLER_11_67 VPWR VGND sg13g2_fill_1
X_07178_ _02952_ net3437 net1009 _00922_ VPWR VGND sg13g2_mux2_1
XFILLER_105_445 VPWR VGND sg13g2_decap_8
X_06129_ net3005 net3014 net1043 _00298_ VPWR VGND sg13g2_mux2_1
XFILLER_106_979 VPWR VGND sg13g2_decap_8
Xclkbuf_4_15_0_clk_regs clknet_0_clk_regs clknet_4_15_0_clk_regs VPWR VGND sg13g2_buf_8
X_08726__1262 VPWR VGND net1682 sg13g2_tiehi
XFILLER_101_684 VPWR VGND sg13g2_decap_4
X_07918__730 VPWR VGND net730 sg13g2_tiehi
X_08621__1355 VPWR VGND net1775 sg13g2_tiehi
XFILLER_46_226 VPWR VGND sg13g2_fill_1
XFILLER_43_933 VPWR VGND sg13g2_fill_2
X_08948__1034 VPWR VGND net1454 sg13g2_tiehi
XFILLER_70_774 VPWR VGND sg13g2_fill_1
XFILLER_42_487 VPWR VGND sg13g2_fill_2
Xinput17 uio_in[7] net17 VPWR VGND sg13g2_buf_2
X_07925__723 VPWR VGND net723 sg13g2_tiehi
XFILLER_7_867 VPWR VGND sg13g2_fill_1
XFILLER_93_866 VPWR VGND sg13g2_fill_2
X_07932__716 VPWR VGND net716 sg13g2_tiehi
X_06480_ net2578 net2081 net1023 _00561_ VPWR VGND sg13g2_mux2_1
X_05500_ net1278 _01386_ _02195_ VPWR VGND sg13g2_nor2_1
X_08245__432 VPWR VGND net432 sg13g2_tiehi
X_05431_ net1232 _02128_ _02134_ _02140_ VPWR VGND sg13g2_nor3_1
XFILLER_21_605 VPWR VGND sg13g2_fill_2
X_08804__1184 VPWR VGND net1604 sg13g2_tiehi
X_08150_ net528 VGND VPWR net2564 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[14\]
+ clknet_leaf_141_clk_regs sg13g2_dfrbpq_1
X_05362_ i_exotiny._2034_\[3\] _00017_ _02084_ VPWR VGND sg13g2_xor2_1
X_07101_ net2694 _02942_ net914 _00855_ VPWR VGND sg13g2_mux2_1
X_08081_ net613 VGND VPWR net2407 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[18\]
+ clknet_leaf_87_clk_regs sg13g2_dfrbpq_1
X_05293_ _02016_ _02017_ _02015_ _02019_ VPWR VGND _02018_ sg13g2_nand4_1
XFILLER_106_209 VPWR VGND sg13g2_decap_8
XFILLER_61_0 VPWR VGND sg13g2_fill_2
X_07032_ _02420_ _02564_ _02934_ VPWR VGND sg13g2_nor2_2
XFILLER_103_916 VPWR VGND sg13g2_decap_8
XFILLER_87_115 VPWR VGND sg13g2_fill_1
X_08983_ net1419 VGND VPWR net1990 i_exotiny._1160_\[4\] clknet_leaf_17_clk_regs sg13g2_dfrbpq_1
XFILLER_102_448 VPWR VGND sg13g2_decap_8
X_08252__425 VPWR VGND net425 sg13g2_tiehi
XFILLER_69_863 VPWR VGND sg13g2_fill_1
X_07934_ net714 VGND VPWR net1925 i_exotiny._1924_\[27\] clknet_leaf_30_clk_regs sg13g2_dfrbpq_1
X_07865_ net2804 net3140 net981 _01332_ VPWR VGND sg13g2_mux2_1
XFILLER_56_535 VPWR VGND sg13g2_fill_2
XFILLER_83_365 VPWR VGND sg13g2_fill_2
X_06816_ net1170 VPWR _02834_ VGND net3655 net1185 sg13g2_o21ai_1
X_07796_ net3323 net2751 net893 _01275_ VPWR VGND sg13g2_mux2_1
X_06747_ VGND VPWR _02773_ _02775_ _02776_ net1135 sg13g2_a21oi_1
X_06678_ _02715_ net1270 _01388_ net1137 VPWR VGND sg13g2_and3_1
X_05629_ net1941 net1065 _02293_ VPWR VGND sg13g2_nor2_1
X_08417_ net268 VGND VPWR net2494 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[16\]
+ clknet_leaf_91_clk_regs sg13g2_dfrbpq_1
XFILLER_51_262 VPWR VGND sg13g2_fill_2
XFILLER_24_487 VPWR VGND sg13g2_fill_1
X_08348_ net330 VGND VPWR _00429_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[18\]
+ clknet_leaf_107_clk_regs sg13g2_dfrbpq_1
XFILLER_20_660 VPWR VGND sg13g2_fill_2
X_08279_ net399 VGND VPWR _00360_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[13\]
+ clknet_leaf_99_clk_regs sg13g2_dfrbpq_1
XFILLER_4_848 VPWR VGND sg13g2_decap_8
X_08437__248 VPWR VGND net248 sg13g2_tiehi
XFILLER_106_776 VPWR VGND sg13g2_decap_8
XFILLER_105_242 VPWR VGND sg13g2_decap_8
Xfanout1104 _02502_ net1104 VPWR VGND sg13g2_buf_1
X_07955__705 VPWR VGND net705 sg13g2_tiehi
Xfanout1126 _01550_ net1126 VPWR VGND sg13g2_buf_8
XFILLER_78_137 VPWR VGND sg13g2_fill_2
Xfanout1115 net1116 net1115 VPWR VGND sg13g2_buf_1
Xfanout1137 _01507_ net1137 VPWR VGND sg13g2_buf_8
Xfanout1159 net1160 net1159 VPWR VGND sg13g2_buf_8
Xfanout1148 _03014_ net1148 VPWR VGND sg13g2_buf_8
XFILLER_47_513 VPWR VGND sg13g2_fill_2
XFILLER_102_993 VPWR VGND sg13g2_decap_8
XFILLER_101_492 VPWR VGND sg13g2_decap_8
XFILLER_93_129 VPWR VGND sg13g2_fill_2
X_08268__410 VPWR VGND net410 sg13g2_tiehi
XFILLER_103_80 VPWR VGND sg13g2_fill_1
XFILLER_16_966 VPWR VGND sg13g2_fill_1
XFILLER_8_68 VPWR VGND sg13g2_fill_1
Xhold609 _00273_ VPWR VGND net2436 sg13g2_dlygate4sd3_1
X_08275__403 VPWR VGND net403 sg13g2_tiehi
XFILLER_98_958 VPWR VGND sg13g2_decap_8
XFILLER_97_457 VPWR VGND sg13g2_fill_1
X_05980_ net2207 net2893 net1048 _00182_ VPWR VGND sg13g2_mux2_1
Xhold1309 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[30\]
+ VPWR VGND net3136 sg13g2_dlygate4sd3_1
X_04931_ _01663_ _01624_ i_exotiny._0040_\[3\] _01619_ i_exotiny._0034_\[3\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_38_546 VPWR VGND sg13g2_fill_1
X_04862_ net3430 VPWR _01596_ VGND net1111 _01583_ sg13g2_o21ai_1
XFILLER_65_354 VPWR VGND sg13g2_fill_1
X_07650_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[23\]
+ net2349 net896 _01158_ VPWR VGND sg13g2_mux2_1
X_07581_ net3627 _03158_ _03159_ VPWR VGND sg13g2_and2_1
X_04793_ _01542_ VPWR _00013_ VGND _01540_ _01541_ sg13g2_o21ai_1
X_06601_ i_exotiny._0314_\[13\] net1160 _02657_ VPWR VGND sg13g2_nor2_1
X_08999__983 VPWR VGND net1403 sg13g2_tiehi
X_06532_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[21\]
+ net2623 net931 _00607_ VPWR VGND sg13g2_mux2_1
X_09251_ net556 VGND VPWR _01306_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[9\]
+ clknet_leaf_128_clk_regs sg13g2_dfrbpq_1
X_06463_ i_exotiny._0039_\[0\] net886 _02608_ _02610_ VPWR VGND sg13g2_mux2_1
X_08202_ net475 VGND VPWR net2318 i_exotiny._0037_\[1\] clknet_leaf_154_clk_regs sg13g2_dfrbpq_2
X_09182_ net799 VGND VPWR _01237_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[4\]
+ clknet_leaf_78_clk_regs sg13g2_dfrbpq_1
X_05414_ VGND VPWR i_exotiny._2034_\[9\] _02123_ _02124_ net1113 sg13g2_a21oi_1
X_06394_ net1071 net3787 _02580_ _00510_ VPWR VGND sg13g2_a21o_1
X_08133_ net1177 VGND VPWR net3544 _00021_ clknet_leaf_48_clk_regs sg13g2_dfrbpq_2
X_05345_ _02068_ _02061_ _02058_ _02069_ VPWR VGND sg13g2_a21o_1
XFILLER_88_1014 VPWR VGND sg13g2_decap_8
X_08064_ net630 VGND VPWR net3030 i_exotiny._0020_\[1\] clknet_leaf_93_clk_regs sg13g2_dfrbpq_2
X_07015_ net2912 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[23\]
+ net918 _00782_ VPWR VGND sg13g2_mux2_1
X_05276_ _02002_ _01790_ i_exotiny._0034_\[0\] _01774_ i_exotiny._0018_\[0\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_102_245 VPWR VGND sg13g2_decap_8
X_08966_ net1436 VGND VPWR _01024_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[2\]
+ clknet_leaf_12_clk_regs sg13g2_dfrbpq_1
Xhold1810 i_exotiny._1160_\[23\] VPWR VGND net3637 sg13g2_dlygate4sd3_1
Xhold1854 i_exotiny.i_rstctl.cnt\[5\] VPWR VGND net3681 sg13g2_dlygate4sd3_1
X_07917_ net731 VGND VPWR net2007 i_exotiny._1924_\[10\] clknet_leaf_33_clk_regs sg13g2_dfrbpq_1
Xhold1832 i_exotiny.i_wb_spi.dat_rx_r\[26\] VPWR VGND net3659 sg13g2_dlygate4sd3_1
X_08897_ net1505 VGND VPWR net3617 i_exotiny.i_wb_spi.dat_rx_r\[27\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_1
Xhold1843 i_exotiny._0315_\[8\] VPWR VGND net3670 sg13g2_dlygate4sd3_1
Xhold1821 _02575_ VPWR VGND net3648 sg13g2_dlygate4sd3_1
Xhold1887 i_exotiny.i_wdg_top.o_wb_dat\[7\] VPWR VGND net3714 sg13g2_dlygate4sd3_1
Xhold1876 i_exotiny.i_wb_spi.cnt_hbit_r\[5\] VPWR VGND net3703 sg13g2_dlygate4sd3_1
X_09290__1399 VPWR VGND net1819 sg13g2_tiehi
XFILLER_17_708 VPWR VGND sg13g2_fill_1
Xhold1865 i_exotiny._0315_\[7\] VPWR VGND net3692 sg13g2_dlygate4sd3_1
X_07848_ net2471 net3134 net987 _01321_ VPWR VGND sg13g2_mux2_1
X_07915__733 VPWR VGND net733 sg13g2_tiehi
Xhold1898 _01113_ VPWR VGND net3725 sg13g2_dlygate4sd3_1
X_07779_ _03213_ net3050 net989 _01262_ VPWR VGND sg13g2_mux2_1
Xclkbuf_leaf_127_clk_regs clknet_5_21__leaf_clk_regs clknet_leaf_127_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_13_969 VPWR VGND sg13g2_decap_8
X_08898__1084 VPWR VGND net1504 sg13g2_tiehi
X_07922__726 VPWR VGND net726 sg13g2_tiehi
XFILLER_4_656 VPWR VGND sg13g2_fill_2
XFILLER_106_573 VPWR VGND sg13g2_decap_8
XFILLER_0_840 VPWR VGND sg13g2_decap_8
X_08235__442 VPWR VGND net442 sg13g2_tiehi
XFILLER_102_790 VPWR VGND sg13g2_decap_8
Xhold6 i_exotiny._2055_\[1\] VPWR VGND net1833 sg13g2_dlygate4sd3_1
XFILLER_48_877 VPWR VGND sg13g2_fill_1
XFILLER_16_752 VPWR VGND sg13g2_fill_2
X_08562__80 VPWR VGND net80 sg13g2_tiehi
XFILLER_31_722 VPWR VGND sg13g2_fill_1
X_08685__1303 VPWR VGND net1723 sg13g2_tiehi
X_08242__435 VPWR VGND net435 sg13g2_tiehi
XFILLER_8_951 VPWR VGND sg13g2_decap_8
X_05130_ _01860_ _01848_ _01859_ VPWR VGND sg13g2_nand2_1
Xhold417 _00733_ VPWR VGND net2244 sg13g2_dlygate4sd3_1
Xhold406 _00531_ VPWR VGND net2233 sg13g2_dlygate4sd3_1
Xhold428 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[6\]
+ VPWR VGND net2255 sg13g2_dlygate4sd3_1
Xhold439 _00712_ VPWR VGND net2266 sg13g2_dlygate4sd3_1
X_05061_ _01793_ _01791_ i_exotiny._0026_\[3\] _01785_ i_exotiny._0043_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_08820_ net1588 VGND VPWR _00878_ i_exotiny.i_wb_spi.state_r\[19\] clknet_leaf_42_clk_regs
+ sg13g2_dfrbpq_1
Xfanout908 net912 net908 VPWR VGND sg13g2_buf_8
Xfanout919 net923 net919 VPWR VGND sg13g2_buf_1
XFILLER_100_705 VPWR VGND sg13g2_fill_1
XFILLER_58_608 VPWR VGND sg13g2_fill_2
Xhold1106 i_exotiny._0038_\[0\] VPWR VGND net2933 sg13g2_dlygate4sd3_1
XFILLER_24_0 VPWR VGND sg13g2_fill_1
X_05963_ i_exotiny._0020_\[0\] net888 _02486_ _02488_ VPWR VGND sg13g2_mux2_1
XFILLER_85_438 VPWR VGND sg13g2_fill_2
X_08751_ net1657 VGND VPWR _00809_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[14\]
+ clknet_leaf_85_clk_regs sg13g2_dfrbpq_1
Xhold1117 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[9\]
+ VPWR VGND net2944 sg13g2_dlygate4sd3_1
Xhold1139 _00612_ VPWR VGND net2966 sg13g2_dlygate4sd3_1
Xhold1128 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[21\]
+ VPWR VGND net2955 sg13g2_dlygate4sd3_1
X_05894_ net1158 VPWR _02479_ VGND _02423_ _02478_ sg13g2_o21ai_1
X_08682_ net1726 VGND VPWR _00740_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[9\]
+ clknet_leaf_116_clk_regs sg13g2_dfrbpq_1
X_04914_ net1255 _01613_ _01640_ _01646_ VPWR VGND sg13g2_nor3_2
X_07702_ VGND VPWR net1142 _03199_ _03200_ net1163 sg13g2_a21oi_1
XFILLER_94_983 VPWR VGND sg13g2_decap_8
X_04845_ net1840 net1111 _01583_ i_exotiny._1902_\[0\] VPWR VGND sg13g2_nor3_1
XFILLER_65_151 VPWR VGND sg13g2_fill_2
X_07633_ net2462 net2686 net897 _01141_ VPWR VGND sg13g2_mux2_1
XFILLER_38_365 VPWR VGND sg13g2_fill_1
XFILLER_0_1022 VPWR VGND sg13g2_decap_8
X_08427__258 VPWR VGND net258 sg13g2_tiehi
X_07564_ net3699 net1231 _03148_ VPWR VGND sg13g2_nor2_1
X_04776_ _01527_ net3724 _01488_ _01490_ VPWR VGND sg13g2_and3_1
XFILLER_41_519 VPWR VGND sg13g2_fill_2
X_09303_ net1357 VGND VPWR net3098 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[29\]
+ clknet_leaf_178_clk_regs sg13g2_dfrbpq_1
X_06515_ net2835 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[8\]
+ net932 _00590_ VPWR VGND sg13g2_mux2_1
X_07495_ net3665 net3670 net902 _01078_ VPWR VGND sg13g2_mux2_1
XFILLER_22_777 VPWR VGND sg13g2_fill_1
X_09234_ net745 VGND VPWR _01289_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[24\]
+ clknet_leaf_135_clk_regs sg13g2_dfrbpq_1
X_06446_ net2206 net2057 net935 _00533_ VPWR VGND sg13g2_mux2_1
X_09165_ net817 VGND VPWR net2749 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[21\]
+ clknet_leaf_174_clk_regs sg13g2_dfrbpq_1
X_06377_ net3343 net879 _02565_ _02569_ VPWR VGND sg13g2_mux2_1
X_08116_ net578 VGND VPWR net2670 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[21\]
+ clknet_leaf_124_clk_regs sg13g2_dfrbpq_1
X_09096_ net1306 VGND VPWR net2786 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[16\]
+ clknet_leaf_142_clk_regs sg13g2_dfrbpq_1
X_05328_ _02052_ _02049_ _02050_ _01979_ _01978_ VPWR VGND sg13g2_a22oi_1
X_08047_ net647 VGND VPWR net2358 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[16\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
Xhold940 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[8\]
+ VPWR VGND net2767 sg13g2_dlygate4sd3_1
X_05259_ _01983_ _01715_ _01701_ _01985_ VPWR VGND sg13g2_a21o_1
Xhold962 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[11\]
+ VPWR VGND net2789 sg13g2_dlygate4sd3_1
Xhold951 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[24\]
+ VPWR VGND net2778 sg13g2_dlygate4sd3_1
Xhold973 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[31\]
+ VPWR VGND net2800 sg13g2_dlygate4sd3_1
XFILLER_103_521 VPWR VGND sg13g2_decap_8
XFILLER_89_755 VPWR VGND sg13g2_fill_2
Xhold995 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[15\]
+ VPWR VGND net2822 sg13g2_dlygate4sd3_1
Xhold984 _01354_ VPWR VGND net2811 sg13g2_dlygate4sd3_1
XFILLER_103_565 VPWR VGND sg13g2_fill_1
X_08949_ net1453 VGND VPWR _01007_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[15\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
Xhold1640 _00696_ VPWR VGND net3467 sg13g2_dlygate4sd3_1
X_08763__1225 VPWR VGND net1645 sg13g2_tiehi
Xhold1651 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[10\]
+ VPWR VGND net3478 sg13g2_dlygate4sd3_1
Xhold1662 i_exotiny._0314_\[21\] VPWR VGND net3489 sg13g2_dlygate4sd3_1
X_08589__1387 VPWR VGND net1807 sg13g2_tiehi
Xhold1684 _00014_ VPWR VGND net3511 sg13g2_dlygate4sd3_1
XFILLER_56_173 VPWR VGND sg13g2_fill_1
Xhold1695 _00007_ VPWR VGND net3522 sg13g2_dlygate4sd3_1
XFILLER_17_516 VPWR VGND sg13g2_decap_8
Xhold1673 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[9\]
+ VPWR VGND net3500 sg13g2_dlygate4sd3_1
XFILLER_32_508 VPWR VGND sg13g2_fill_1
XFILLER_44_42 VPWR VGND sg13g2_decap_4
XFILLER_12_210 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_95_clk_regs clknet_5_28__leaf_clk_regs clknet_leaf_95_clk_regs VPWR VGND
+ sg13g2_buf_8
Xclkbuf_leaf_24_clk_regs clknet_5_12__leaf_clk_regs clknet_leaf_24_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_5_910 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_fill_2
XFILLER_5_987 VPWR VGND sg13g2_decap_8
X_08989__993 VPWR VGND net1413 sg13g2_tiehi
XFILLER_106_370 VPWR VGND sg13g2_decap_8
X_08272__406 VPWR VGND net406 sg13g2_tiehi
XFILLER_67_438 VPWR VGND sg13g2_fill_1
XFILLER_91_931 VPWR VGND sg13g2_decap_8
XFILLER_63_611 VPWR VGND sg13g2_fill_2
XFILLER_63_600 VPWR VGND sg13g2_fill_1
X_04630_ VPWR _01392_ net3788 VGND sg13g2_inv_1
XFILLER_50_349 VPWR VGND sg13g2_fill_1
X_08996__986 VPWR VGND net1406 sg13g2_tiehi
X_07280_ net2654 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[9\]
+ net908 _00997_ VPWR VGND sg13g2_mux2_1
X_06300_ net3274 net878 _02552_ _02556_ VPWR VGND sg13g2_mux2_1
XFILLER_31_563 VPWR VGND sg13g2_fill_1
X_06231_ net3515 i_exotiny._0031_\[1\] net1040 _00380_ VPWR VGND sg13g2_mux2_1
XFILLER_102_1000 VPWR VGND sg13g2_decap_8
X_06162_ net2557 net3149 net952 _00324_ VPWR VGND sg13g2_mux2_1
Xhold203 _01122_ VPWR VGND net2030 sg13g2_dlygate4sd3_1
XFILLER_85_1006 VPWR VGND sg13g2_decap_8
X_06093_ net2073 net2855 net960 _00269_ VPWR VGND sg13g2_mux2_1
Xhold225 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[22\]
+ VPWR VGND net2052 sg13g2_dlygate4sd3_1
Xhold214 _01051_ VPWR VGND net2041 sg13g2_dlygate4sd3_1
X_05113_ _01385_ VPWR _01843_ VGND _01841_ _01842_ sg13g2_o21ai_1
Xhold269 _00379_ VPWR VGND net2096 sg13g2_dlygate4sd3_1
Xhold236 i_exotiny._1614_\[0\] VPWR VGND net2063 sg13g2_dlygate4sd3_1
Xhold247 _00265_ VPWR VGND net2074 sg13g2_dlygate4sd3_1
Xhold258 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[8\]
+ VPWR VGND net2085 sg13g2_dlygate4sd3_1
X_05044_ _01756_ _01768_ _01776_ VPWR VGND sg13g2_nor2_2
XFILLER_98_563 VPWR VGND sg13g2_fill_2
X_08803_ net1605 VGND VPWR _00861_ i_exotiny.i_wb_spi.state_r\[2\] clknet_leaf_44_clk_regs
+ sg13g2_dfrbpq_1
X_08734_ net1674 VGND VPWR _00792_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[29\]
+ clknet_leaf_121_clk_regs sg13g2_dfrbpq_1
X_06995_ _02928_ net1141 net1165 _02929_ VPWR VGND sg13g2_a21o_1
X_05946_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[11\]
+ net2822 net969 _00155_ VPWR VGND sg13g2_mux2_1
X_08665_ net1203 VGND VPWR i_exotiny._2043_\[2\] i_exotiny._2034_\[2\] net1228 sg13g2_dfrbpq_2
X_05877_ net3282 net876 _02421_ _02464_ VPWR VGND sg13g2_mux2_1
X_04828_ net1863 net1851 net1861 net1848 _01568_ VPWR VGND sg13g2_nor4_1
X_07616_ net2054 _03180_ _03181_ VPWR VGND sg13g2_nor2_1
X_08596_ net1800 VGND VPWR net3809 i_exotiny._1612_\[0\] clknet_leaf_24_clk_regs sg13g2_dfrbpq_2
X_07912__736 VPWR VGND net736 sg13g2_tiehi
X_07547_ _03137_ net1883 net3586 net2298 VPWR VGND sg13g2_and3_1
X_04759_ _01509_ net1218 _01487_ _01510_ VPWR VGND sg13g2_a21o_2
XFILLER_41_338 VPWR VGND sg13g2_fill_1
X_07478_ _03105_ net3819 _03104_ VPWR VGND sg13g2_nand2_1
X_06429_ net1146 _02593_ net1219 _02606_ VPWR VGND sg13g2_nand3_1
X_08225__452 VPWR VGND net452 sg13g2_tiehi
X_09217_ net762 VGND VPWR net3293 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[7\]
+ clknet_leaf_134_clk_regs sg13g2_dfrbpq_1
X_09148_ net834 VGND VPWR net2991 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[4\]
+ clknet_leaf_174_clk_regs sg13g2_dfrbpq_1
XFILLER_5_217 VPWR VGND sg13g2_fill_1
X_09079_ net1323 VGND VPWR _01134_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[19\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_08817__1171 VPWR VGND net1591 sg13g2_tiehi
Xhold770 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[15\]
+ VPWR VGND net2597 sg13g2_dlygate4sd3_1
Xhold781 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[26\]
+ VPWR VGND net2608 sg13g2_dlygate4sd3_1
XFILLER_2_957 VPWR VGND sg13g2_decap_8
XFILLER_104_874 VPWR VGND sg13g2_decap_8
Xhold792 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[18\]
+ VPWR VGND net2619 sg13g2_dlygate4sd3_1
XFILLER_7_1017 VPWR VGND sg13g2_decap_8
XFILLER_103_395 VPWR VGND sg13g2_decap_8
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
XFILLER_76_257 VPWR VGND sg13g2_fill_1
X_08232__445 VPWR VGND net445 sg13g2_tiehi
Xclkbuf_leaf_142_clk_regs clknet_5_17__leaf_clk_regs clknet_leaf_142_clk_regs VPWR
+ VGND sg13g2_buf_8
Xhold1470 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[8\]
+ VPWR VGND net3297 sg13g2_dlygate4sd3_1
XFILLER_17_313 VPWR VGND sg13g2_fill_2
XFILLER_45_600 VPWR VGND sg13g2_fill_1
Xhold1492 i_exotiny._0030_\[1\] VPWR VGND net3319 sg13g2_dlygate4sd3_1
Xhold1481 i_exotiny._1611_\[18\] VPWR VGND net3308 sg13g2_dlygate4sd3_1
XFILLER_45_633 VPWR VGND sg13g2_fill_2
X_08087__607 VPWR VGND net607 sg13g2_tiehi
XFILLER_73_986 VPWR VGND sg13g2_fill_2
XFILLER_44_132 VPWR VGND sg13g2_fill_1
XFILLER_45_699 VPWR VGND sg13g2_decap_4
XFILLER_41_861 VPWR VGND sg13g2_fill_1
XFILLER_9_545 VPWR VGND sg13g2_fill_1
X_08417__268 VPWR VGND net268 sg13g2_tiehi
XFILLER_95_511 VPWR VGND sg13g2_fill_2
X_05800_ _01473_ _01683_ _01467_ _02417_ VPWR VGND _02416_ sg13g2_nand4_1
X_06780_ VGND VPWR net2012 net1131 _02804_ _02803_ sg13g2_a21oi_1
X_05731_ _02369_ net1972 net1073 VPWR VGND sg13g2_nand2_1
X_05662_ VGND VPWR net1063 _02317_ _00041_ _02315_ sg13g2_a21oi_1
X_08450_ net230 VGND VPWR _00524_ i_exotiny._0039_\[2\] clknet_leaf_114_clk_regs sg13g2_dfrbpq_2
X_04613_ VPWR _01375_ _00016_ VGND sg13g2_inv_1
X_08381_ net297 VGND VPWR net2001 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[19\]
+ clknet_leaf_134_clk_regs sg13g2_dfrbpq_1
X_07401_ VGND VPWR i_exotiny._0369_\[12\] net1147 _03053_ _03052_ sg13g2_a21oi_1
XFILLER_51_669 VPWR VGND sg13g2_decap_8
X_05593_ _01978_ VPWR _02267_ VGND _01980_ _02266_ sg13g2_o21ai_1
X_07332_ VGND VPWR i_exotiny._0369_\[5\] _02994_ _02996_ i_exotiny._0369_\[20\] sg13g2_a21oi_1
X_07263_ net2614 net2973 net1003 _00986_ VPWR VGND sg13g2_mux2_1
X_06214_ net2774 net3427 net945 _00369_ VPWR VGND sg13g2_mux2_1
X_07194_ net3576 net3574 net1093 _00930_ VPWR VGND sg13g2_mux2_1
X_09002_ net1400 VGND VPWR _01060_ i_exotiny._1160_\[23\] clknet_leaf_161_clk_regs
+ sg13g2_dfrbpq_1
X_06145_ i_exotiny._0037_\[2\] net877 _02526_ _02530_ VPWR VGND sg13g2_mux2_1
X_06076_ i_exotiny._0038_\[2\] net2255 net959 _00252_ VPWR VGND sg13g2_mux2_1
XFILLER_104_159 VPWR VGND sg13g2_decap_8
X_05027_ _01759_ i_exotiny._0079_\[3\] VPWR VGND i_exotiny._0079_\[2\] sg13g2_nand2b_2
XFILLER_101_822 VPWR VGND sg13g2_decap_8
XFILLER_100_332 VPWR VGND sg13g2_decap_8
XFILLER_101_899 VPWR VGND sg13g2_decap_8
X_06978_ net2908 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[24\]
+ net1021 _00751_ VPWR VGND sg13g2_mux2_1
X_05929_ net872 i_exotiny._0019_\[3\] _02478_ _02483_ VPWR VGND sg13g2_mux2_1
X_08717_ net1691 VGND VPWR _00775_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[12\]
+ clknet_leaf_119_clk_regs sg13g2_dfrbpq_1
X_08648_ net1749 VGND VPWR _00716_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[17\]
+ clknet_leaf_148_clk_regs sg13g2_dfrbpq_1
XFILLER_15_806 VPWR VGND sg13g2_fill_2
XFILLER_42_636 VPWR VGND sg13g2_fill_1
XFILLER_42_647 VPWR VGND sg13g2_decap_4
X_08579_ net1824 VGND VPWR _00652_ i_exotiny._0314_\[24\] clknet_leaf_0_clk_regs sg13g2_dfrbpq_1
XFILLER_14_349 VPWR VGND sg13g2_fill_1
XFILLER_41_179 VPWR VGND sg13g2_fill_2
XFILLER_50_691 VPWR VGND sg13g2_decap_8
XFILLER_96_308 VPWR VGND sg13g2_decap_8
XFILLER_2_754 VPWR VGND sg13g2_decap_8
X_08986__996 VPWR VGND net1416 sg13g2_tiehi
XFILLER_104_682 VPWR VGND sg13g2_fill_1
XFILLER_104_671 VPWR VGND sg13g2_decap_8
XFILLER_103_192 VPWR VGND sg13g2_decap_8
XFILLER_45_430 VPWR VGND sg13g2_fill_2
X_08840__1146 VPWR VGND net1566 sg13g2_tiehi
XFILLER_33_603 VPWR VGND sg13g2_fill_2
XFILLER_33_625 VPWR VGND sg13g2_decap_4
XFILLER_14_883 VPWR VGND sg13g2_fill_1
X_08993__989 VPWR VGND net1409 sg13g2_tiehi
XFILLER_9_353 VPWR VGND sg13g2_fill_2
X_07950_ net706 VGND VPWR net3704 i_exotiny.i_wb_spi.cnt_hbit_r\[5\] clknet_leaf_38_clk_regs
+ sg13g2_dfrbpq_2
X_06901_ _02902_ net1970 net3766 VPWR VGND sg13g2_nand2b_1
X_07881_ net2558 net2938 net980 _01348_ VPWR VGND sg13g2_mux2_1
XFILLER_96_886 VPWR VGND sg13g2_decap_8
XFILLER_95_363 VPWR VGND sg13g2_fill_2
X_06832_ VGND VPWR net1096 _02846_ _00681_ _02847_ sg13g2_a21oi_1
X_08215__462 VPWR VGND net462 sg13g2_tiehi
X_06763_ VGND VPWR _01413_ net1190 _02789_ net1169 sg13g2_a21oi_1
X_08791__1197 VPWR VGND net1617 sg13g2_tiehi
X_08502_ net178 VGND VPWR _00576_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[22\]
+ clknet_leaf_84_clk_regs sg13g2_dfrbpq_1
X_05714_ VGND VPWR net1059 _02355_ _00054_ _02356_ sg13g2_a21oi_1
X_09098__884 VPWR VGND net1304 sg13g2_tiehi
XFILLER_63_282 VPWR VGND sg13g2_fill_2
X_08980__1002 VPWR VGND net1422 sg13g2_tiehi
X_06694_ net3632 net1102 _02731_ VPWR VGND sg13g2_nor2_1
X_05645_ VGND VPWR i_exotiny._1615_\[3\] net1124 _02305_ _02304_ sg13g2_a21oi_1
XFILLER_12_809 VPWR VGND sg13g2_fill_2
X_08433_ net252 VGND VPWR _00507_ i_exotiny._0369_\[24\] clknet_leaf_16_clk_regs sg13g2_dfrbpq_1
X_08364_ net314 VGND VPWR _00445_ i_exotiny._0014_\[2\] clknet_leaf_140_clk_regs sg13g2_dfrbpq_2
X_05576_ i_exotiny._1489_\[2\] net1985 _02255_ _02253_ _01385_ VPWR VGND sg13g2_a22oi_1
X_07315_ net1249 net3800 net1150 _01027_ VPWR VGND sg13g2_mux2_1
X_08295_ net383 VGND VPWR _00376_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[29\]
+ clknet_leaf_106_clk_regs sg13g2_dfrbpq_1
X_07246_ net3089 net2934 net1005 _00969_ VPWR VGND sg13g2_mux2_1
X_08222__455 VPWR VGND net455 sg13g2_tiehi
X_07177_ i_exotiny._0036_\[3\] net872 _02947_ _02952_ VPWR VGND sg13g2_mux2_1
XFILLER_106_958 VPWR VGND sg13g2_decap_8
XFILLER_105_424 VPWR VGND sg13g2_decap_8
X_08077__617 VPWR VGND net617 sg13g2_tiehi
X_06128_ net3454 net2602 net1044 _00297_ VPWR VGND sg13g2_mux2_1
X_06059_ net2800 net2657 net963 _00244_ VPWR VGND sg13g2_mux2_1
XFILLER_59_555 VPWR VGND sg13g2_fill_2
XFILLER_4_1009 VPWR VGND sg13g2_decap_8
XFILLER_46_238 VPWR VGND sg13g2_fill_2
XFILLER_27_441 VPWR VGND sg13g2_fill_1
XFILLER_55_794 VPWR VGND sg13g2_fill_2
XFILLER_36_98 VPWR VGND sg13g2_fill_2
X_08407__278 VPWR VGND net278 sg13g2_tiehi
XFILLER_70_797 VPWR VGND sg13g2_fill_2
XFILLER_35_1000 VPWR VGND sg13g2_fill_2
X_08858__1128 VPWR VGND net1548 sg13g2_tiehi
XFILLER_96_127 VPWR VGND sg13g2_fill_2
XFILLER_2_584 VPWR VGND sg13g2_fill_1
XFILLER_78_853 VPWR VGND sg13g2_fill_1
XFILLER_28_7 VPWR VGND sg13g2_fill_2
XFILLER_37_216 VPWR VGND sg13g2_fill_1
XFILLER_93_878 VPWR VGND sg13g2_fill_2
XFILLER_80_528 VPWR VGND sg13g2_fill_2
X_05430_ VGND VPWR i_exotiny._1615_\[0\] _02136_ _02139_ _02137_ sg13g2_a21oi_1
X_08776__1212 VPWR VGND net1632 sg13g2_tiehi
X_05361_ i_exotiny._2034_\[5\] _00019_ _02083_ VPWR VGND sg13g2_xor2_1
X_07100_ net3063 net886 _02940_ _02942_ VPWR VGND sg13g2_mux2_1
X_08080_ net614 VGND VPWR _00161_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[17\]
+ clknet_leaf_91_clk_regs sg13g2_dfrbpq_1
X_05292_ _02018_ _01634_ i_exotiny._0013_\[0\] _01627_ i_exotiny._0028_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_07031_ net3301 _02933_ net919 _00794_ VPWR VGND sg13g2_mux2_1
XFILLER_102_427 VPWR VGND sg13g2_decap_8
X_08982_ net1420 VGND VPWR net1950 i_exotiny._1160_\[3\] clknet_leaf_15_clk_regs sg13g2_dfrbpq_1
X_07933_ net715 VGND VPWR net1983 i_exotiny._1924_\[26\] clknet_leaf_30_clk_regs sg13g2_dfrbpq_1
X_07864_ i_exotiny._0021_\[2\] net2451 net981 _01331_ VPWR VGND sg13g2_mux2_1
XFILLER_28_205 VPWR VGND sg13g2_fill_2
XFILLER_96_694 VPWR VGND sg13g2_fill_2
XFILLER_83_322 VPWR VGND sg13g2_fill_2
XFILLER_56_525 VPWR VGND sg13g2_fill_1
X_06815_ net3505 net1189 _02833_ VPWR VGND sg13g2_nor2_1
X_07795_ net2833 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[13\]
+ net894 _01274_ VPWR VGND sg13g2_mux2_1
X_06746_ _02774_ VPWR _02775_ VGND net3778 net1190 sg13g2_o21ai_1
X_06677_ VGND VPWR _01362_ _02712_ _02714_ _02713_ sg13g2_a21oi_1
X_08416_ net269 VGND VPWR net2852 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[15\]
+ clknet_leaf_97_clk_regs sg13g2_dfrbpq_1
X_05628_ VGND VPWR i_exotiny._1612_\[3\] net1124 _02292_ _02291_ sg13g2_a21oi_1
XFILLER_52_764 VPWR VGND sg13g2_fill_1
XFILLER_40_915 VPWR VGND sg13g2_fill_1
XFILLER_40_926 VPWR VGND sg13g2_fill_2
X_08347_ net331 VGND VPWR _00428_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[17\]
+ clknet_leaf_94_clk_regs sg13g2_dfrbpq_1
X_05559_ _02241_ net3729 net1071 VPWR VGND sg13g2_nand2_1
X_08278_ net400 VGND VPWR _00359_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[12\]
+ clknet_leaf_101_clk_regs sg13g2_dfrbpq_1
XFILLER_22_45 VPWR VGND sg13g2_fill_2
X_07229_ i_exotiny.i_wb_spi.dat_rx_r\[25\] net3659 net1086 _00954_ VPWR VGND sg13g2_mux2_1
X_08639__1338 VPWR VGND net1758 sg13g2_tiehi
XFILLER_4_827 VPWR VGND sg13g2_decap_8
XFILLER_106_755 VPWR VGND sg13g2_decap_8
XFILLER_105_221 VPWR VGND sg13g2_decap_8
XFILLER_65_1026 VPWR VGND sg13g2_fill_2
XFILLER_79_617 VPWR VGND sg13g2_fill_1
XFILLER_105_298 VPWR VGND sg13g2_decap_8
Xfanout1127 _00026_ net1127 VPWR VGND sg13g2_buf_8
Xfanout1105 i_exotiny._2160_ net1105 VPWR VGND sg13g2_buf_8
Xfanout1116 net1117 net1116 VPWR VGND sg13g2_buf_8
Xfanout1138 net1141 net1138 VPWR VGND sg13g2_buf_8
XFILLER_102_972 VPWR VGND sg13g2_decap_8
Xfanout1149 _03014_ net1149 VPWR VGND sg13g2_buf_1
X_08983__999 VPWR VGND net1419 sg13g2_tiehi
XFILLER_101_471 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_49_clk_regs clknet_5_14__leaf_clk_regs clknet_leaf_49_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_43_720 VPWR VGND sg13g2_decap_4
XFILLER_63_52 VPWR VGND sg13g2_fill_2
XFILLER_43_764 VPWR VGND sg13g2_fill_1
XFILLER_70_594 VPWR VGND sg13g2_fill_1
XFILLER_7_621 VPWR VGND sg13g2_fill_1
XFILLER_6_153 VPWR VGND sg13g2_fill_1
X_08205__472 VPWR VGND net472 sg13g2_tiehi
XFILLER_6_164 VPWR VGND sg13g2_fill_1
X_09088__894 VPWR VGND net1314 sg13g2_tiehi
XFILLER_98_937 VPWR VGND sg13g2_decap_8
XFILLER_97_436 VPWR VGND sg13g2_decap_8
XFILLER_69_127 VPWR VGND sg13g2_fill_2
XFILLER_3_893 VPWR VGND sg13g2_decap_8
X_04930_ _01657_ _01660_ _01635_ _01662_ VPWR VGND _01661_ sg13g2_nand4_1
XFILLER_93_675 VPWR VGND sg13g2_fill_2
X_04861_ _01595_ _01579_ _01594_ _01575_ i_exotiny.i_wb_spi.cnt_presc_r\[6\] VPWR
+ VGND sg13g2_a22oi_1
X_07580_ net1204 net1886 _03158_ _01118_ VPWR VGND sg13g2_nor3_1
X_06600_ net1194 _02655_ _02656_ _00640_ VPWR VGND sg13g2_nor3_1
X_08212__465 VPWR VGND net465 sg13g2_tiehi
X_04792_ net3702 _01487_ net1281 _01542_ VPWR VGND sg13g2_nand3_1
X_06531_ net2701 net2919 net933 _00606_ VPWR VGND sg13g2_mux2_1
X_08067__627 VPWR VGND net627 sg13g2_tiehi
X_09095__887 VPWR VGND net1307 sg13g2_tiehi
X_09250_ net557 VGND VPWR _01305_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[8\]
+ clknet_leaf_126_clk_regs sg13g2_dfrbpq_1
X_08201_ net476 VGND VPWR net3112 i_exotiny._0037_\[0\] clknet_leaf_151_clk_regs sg13g2_dfrbpq_2
X_06462_ net3346 net3115 net935 _00549_ VPWR VGND sg13g2_mux2_1
X_09181_ net800 VGND VPWR _01236_ i_exotiny._0026_\[3\] clknet_leaf_76_clk_regs sg13g2_dfrbpq_2
X_05413_ net1113 _02122_ _02123_ i_exotiny._2043_\[8\] VPWR VGND sg13g2_nor3_1
XFILLER_21_447 VPWR VGND sg13g2_fill_1
X_06393_ _02219_ _02572_ _02579_ _02580_ VPWR VGND sg13g2_nor3_1
X_08132_ net1175 VGND VPWR _00213_ _00020_ clknet_leaf_36_clk_regs sg13g2_dfrbpq_2
X_05344_ VPWR VGND _01837_ _02066_ _02067_ _01834_ _02068_ _02065_ sg13g2_a221oi_1
X_08063_ net631 VGND VPWR net2676 i_exotiny._0020_\[0\] clknet_leaf_89_clk_regs sg13g2_dfrbpq_2
X_05275_ _02001_ _01789_ i_exotiny._0024_\[0\] _01765_ i_exotiny._0027_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_07014_ net3093 net3287 net920 _00781_ VPWR VGND sg13g2_mux2_1
XFILLER_89_937 VPWR VGND sg13g2_fill_1
XFILLER_88_425 VPWR VGND sg13g2_fill_2
XFILLER_0_307 VPWR VGND sg13g2_fill_2
XFILLER_103_769 VPWR VGND sg13g2_decap_8
XFILLER_102_224 VPWR VGND sg13g2_decap_8
X_08965_ net1437 VGND VPWR _01023_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[31\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
Xhold1800 i_exotiny.i_wdg_top.clk_div_inst.cnt\[4\] VPWR VGND net3627 sg13g2_dlygate4sd3_1
X_07916_ net732 VGND VPWR net1944 i_exotiny._1924_\[9\] clknet_leaf_33_clk_regs sg13g2_dfrbpq_1
Xhold1811 i_exotiny.i_wb_spi.dat_rx_r\[23\] VPWR VGND net3638 sg13g2_dlygate4sd3_1
Xhold1822 i_exotiny.i_wdg_top.clk_div_inst.cnt\[15\] VPWR VGND net3649 sg13g2_dlygate4sd3_1
Xhold1844 i_exotiny.i_wdg_top.clk_div_inst.cnt\[5\] VPWR VGND net3671 sg13g2_dlygate4sd3_1
Xhold1833 _00954_ VPWR VGND net3660 sg13g2_dlygate4sd3_1
X_08896_ net1506 VGND VPWR net3660 i_exotiny.i_wb_spi.dat_rx_r\[26\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_1
Xhold1855 _02903_ VPWR VGND net3682 sg13g2_dlygate4sd3_1
Xhold1877 _00060_ VPWR VGND net3704 sg13g2_dlygate4sd3_1
XFILLER_17_12 VPWR VGND sg13g2_fill_1
Xhold1866 _01077_ VPWR VGND net3693 sg13g2_dlygate4sd3_1
X_07847_ net2536 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[23\]
+ net983 _01320_ VPWR VGND sg13g2_mux2_1
X_07778_ i_exotiny._0026_\[1\] net883 _03210_ _03213_ VPWR VGND sg13g2_mux2_1
Xhold1888 _02405_ VPWR VGND net3715 sg13g2_dlygate4sd3_1
Xhold1899 i_exotiny._0571_ VPWR VGND net3726 sg13g2_dlygate4sd3_1
XFILLER_71_358 VPWR VGND sg13g2_fill_1
X_06729_ VPWR VGND _01506_ _02757_ _02760_ _01366_ _00665_ net1068 sg13g2_a221oi_1
XFILLER_40_712 VPWR VGND sg13g2_fill_2
XFILLER_12_436 VPWR VGND sg13g2_fill_2
XFILLER_40_734 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_167_clk_regs clknet_5_4__leaf_clk_regs clknet_leaf_167_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_106_552 VPWR VGND sg13g2_decap_8
Xhold7 i_exotiny.i_wb_spi.state_r\[26\] VPWR VGND net1834 sg13g2_dlygate4sd3_1
XFILLER_0_896 VPWR VGND sg13g2_decap_8
XFILLER_75_642 VPWR VGND sg13g2_fill_2
XFILLER_15_285 VPWR VGND sg13g2_fill_1
XFILLER_8_930 VPWR VGND sg13g2_decap_8
XFILLER_12_981 VPWR VGND sg13g2_decap_8
XFILLER_11_480 VPWR VGND sg13g2_fill_1
Xhold407 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[24\]
+ VPWR VGND net2234 sg13g2_dlygate4sd3_1
Xhold418 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[20\]
+ VPWR VGND net2245 sg13g2_dlygate4sd3_1
XFILLER_99_81 VPWR VGND sg13g2_fill_2
Xhold429 _00252_ VPWR VGND net2256 sg13g2_dlygate4sd3_1
X_05060_ net1239 net1241 net1237 _01792_ VGND VPWR _01757_ sg13g2_nor4_2
Xfanout909 net912 net909 VPWR VGND sg13g2_buf_8
X_08750_ net1658 VGND VPWR _00808_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[13\]
+ clknet_5_30__leaf_clk_regs sg13g2_dfrbpq_1
X_05962_ net2726 net2505 net966 _00171_ VPWR VGND sg13g2_mux2_1
Xhold1107 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[9\]
+ VPWR VGND net2934 sg13g2_dlygate4sd3_1
Xhold1118 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[23\]
+ VPWR VGND net2945 sg13g2_dlygate4sd3_1
Xhold1129 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[27\]
+ VPWR VGND net2956 sg13g2_dlygate4sd3_1
XFILLER_94_962 VPWR VGND sg13g2_decap_8
X_05893_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[4\] _02476_ _02478_
+ VPWR VGND i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[3\] sg13g2_nand3b_1
X_08681_ net1727 VGND VPWR net3100 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[8\]
+ clknet_leaf_102_clk_regs sg13g2_dfrbpq_1
X_07701_ _02419_ _02477_ _03199_ VPWR VGND sg13g2_nor2_2
X_04913_ net1222 _01620_ _01623_ _01645_ VPWR VGND sg13g2_nor3_2
X_04844_ net1111 _01583_ _01584_ VPWR VGND sg13g2_nor2_1
XFILLER_0_1001 VPWR VGND sg13g2_decap_8
X_07632_ net2186 net2607 net898 _01140_ VPWR VGND sg13g2_mux2_1
XFILLER_80_122 VPWR VGND sg13g2_fill_2
X_04775_ _01526_ net1283 _01525_ VPWR VGND sg13g2_nand2_1
X_07563_ net3520 _01527_ _02177_ _03146_ _03147_ VPWR VGND sg13g2_nor4_1
X_09302_ net1533 VGND VPWR _01357_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[28\]
+ clknet_leaf_178_clk_regs sg13g2_dfrbpq_1
XFILLER_34_561 VPWR VGND sg13g2_fill_1
X_06514_ i_exotiny._0043_\[3\] net2274 net931 _00589_ VPWR VGND sg13g2_mux2_1
X_07494_ net3626 net3692 net907 _01077_ VPWR VGND sg13g2_mux2_1
X_06445_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[14\]
+ net2550 _02609_ _00532_ VPWR VGND sg13g2_mux2_1
X_09233_ net746 VGND VPWR _01288_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[23\]
+ clknet_leaf_134_clk_regs sg13g2_dfrbpq_1
X_09164_ net818 VGND VPWR net2049 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[20\]
+ clknet_leaf_176_clk_regs sg13g2_dfrbpq_1
X_06376_ _02568_ net2576 net1029 _00504_ VPWR VGND sg13g2_mux2_1
X_08115_ net579 VGND VPWR _00196_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[20\]
+ clknet_leaf_101_clk_regs sg13g2_dfrbpq_1
X_08853__1133 VPWR VGND net1553 sg13g2_tiehi
X_09095_ net1307 VGND VPWR _01150_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[15\]
+ clknet_leaf_144_clk_regs sg13g2_dfrbpq_1
X_05327_ _02049_ _02050_ _02051_ VPWR VGND sg13g2_and2_1
X_08046_ net648 VGND VPWR _00127_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[15\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
Xhold930 _00280_ VPWR VGND net2757 sg13g2_dlygate4sd3_1
X_05258_ VGND VPWR _01371_ _01739_ _01984_ _01983_ sg13g2_a21oi_1
XFILLER_103_500 VPWR VGND sg13g2_decap_8
Xhold963 _01003_ VPWR VGND net2790 sg13g2_dlygate4sd3_1
Xhold941 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[28\]
+ VPWR VGND net2768 sg13g2_dlygate4sd3_1
Xhold952 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[31\]
+ VPWR VGND net2779 sg13g2_dlygate4sd3_1
X_05189_ _01915_ _01736_ _01701_ _01917_ VPWR VGND sg13g2_a21o_1
Xhold985 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[28\]
+ VPWR VGND net2812 sg13g2_dlygate4sd3_1
Xhold996 _00155_ VPWR VGND net2823 sg13g2_dlygate4sd3_1
Xhold974 _00248_ VPWR VGND net2801 sg13g2_dlygate4sd3_1
X_08948_ net1454 VGND VPWR net2036 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[14\]
+ clknet_leaf_75_clk_regs sg13g2_dfrbpq_1
Xhold1641 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[25\]
+ VPWR VGND net3468 sg13g2_dlygate4sd3_1
X_08879_ net1523 VGND VPWR net1934 i_exotiny.i_wb_spi.dat_rx_r\[9\] clknet_leaf_59_clk_regs
+ sg13g2_dfrbpq_1
Xhold1652 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[15\]
+ VPWR VGND net3479 sg13g2_dlygate4sd3_1
Xhold1630 i_exotiny._0369_\[30\] VPWR VGND net3457 sg13g2_dlygate4sd3_1
Xhold1685 _00025_ VPWR VGND net3512 sg13g2_dlygate4sd3_1
Xhold1674 i_exotiny._1616_\[0\] VPWR VGND net3501 sg13g2_dlygate4sd3_1
Xhold1663 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[7\]
+ VPWR VGND net3490 sg13g2_dlygate4sd3_1
Xhold1696 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[0\] VPWR
+ VGND net3523 sg13g2_dlygate4sd3_1
XFILLER_44_325 VPWR VGND sg13g2_fill_1
XFILLER_44_32 VPWR VGND sg13g2_fill_1
XFILLER_9_727 VPWR VGND sg13g2_fill_2
XFILLER_100_60 VPWR VGND sg13g2_fill_1
XFILLER_5_966 VPWR VGND sg13g2_decap_8
X_08202__475 VPWR VGND net475 sg13g2_tiehi
Xclkbuf_leaf_64_clk_regs clknet_5_13__leaf_clk_regs clknet_leaf_64_clk_regs VPWR VGND
+ sg13g2_buf_8
X_09085__897 VPWR VGND net1317 sg13g2_tiehi
X_08057__637 VPWR VGND net637 sg13g2_tiehi
XFILLER_79_266 VPWR VGND sg13g2_fill_1
XFILLER_76_984 VPWR VGND sg13g2_fill_2
XFILLER_36_815 VPWR VGND sg13g2_fill_2
XFILLER_47_174 VPWR VGND sg13g2_fill_2
XFILLER_91_987 VPWR VGND sg13g2_decap_8
XFILLER_90_497 VPWR VGND sg13g2_fill_1
XFILLER_44_881 VPWR VGND sg13g2_fill_2
X_08634__1343 VPWR VGND net1763 sg13g2_tiehi
X_06230_ net2095 i_exotiny._0031_\[0\] net1040 _00379_ VPWR VGND sg13g2_mux2_1
X_06161_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[9\]
+ net2218 net953 _00323_ VPWR VGND sg13g2_mux2_1
X_06092_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[18\]
+ net2413 net958 _00268_ VPWR VGND sg13g2_mux2_1
Xhold215 i_exotiny._1615_\[0\] VPWR VGND net2042 sg13g2_dlygate4sd3_1
Xhold204 i_exotiny._1924_\[17\] VPWR VGND net2031 sg13g2_dlygate4sd3_1
Xhold226 _00909_ VPWR VGND net2053 sg13g2_dlygate4sd3_1
X_05112_ _01840_ _01720_ _01701_ _01842_ VPWR VGND sg13g2_a21o_1
Xhold237 _00215_ VPWR VGND net2064 sg13g2_dlygate4sd3_1
Xhold259 _00084_ VPWR VGND net2086 sg13g2_dlygate4sd3_1
Xhold248 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[17\]
+ VPWR VGND net2075 sg13g2_dlygate4sd3_1
X_05043_ _01775_ i_exotiny._0018_\[3\] _01774_ VPWR VGND sg13g2_nand2_1
X_08433__252 VPWR VGND net252 sg13g2_tiehi
XFILLER_100_514 VPWR VGND sg13g2_decap_8
X_08802_ net1606 VGND VPWR _00860_ i_exotiny.i_wb_spi.state_r\[1\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_58_439 VPWR VGND sg13g2_fill_1
X_06994_ _02517_ _02532_ _02928_ VPWR VGND sg13g2_nor2_2
X_05945_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[10\]
+ net2969 net967 _00154_ VPWR VGND sg13g2_mux2_1
XFILLER_86_759 VPWR VGND sg13g2_fill_1
X_08733_ net1675 VGND VPWR _00791_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[28\]
+ clknet_leaf_117_clk_regs sg13g2_dfrbpq_1
X_08664_ net1203 VGND VPWR i_exotiny._2043_\[1\] i_exotiny._2034_\[1\] net1228 sg13g2_dfrbpq_2
XFILLER_82_954 VPWR VGND sg13g2_fill_1
XFILLER_54_634 VPWR VGND sg13g2_fill_2
X_05876_ _01470_ _02462_ _02463_ VPWR VGND sg13g2_nor2b_2
XFILLER_27_848 VPWR VGND sg13g2_fill_2
X_07615_ net1205 net1881 _03180_ _01131_ VPWR VGND sg13g2_nor3_1
X_04827_ net1869 net1857 net1855 net1847 _01567_ VPWR VGND sg13g2_nor4_1
X_08595_ net1801 VGND VPWR _00667_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data[0]
+ clknet_leaf_24_clk_regs sg13g2_dfrbpq_2
XFILLER_54_667 VPWR VGND sg13g2_fill_1
XFILLER_14_509 VPWR VGND sg13g2_fill_2
X_07546_ VGND VPWR net1883 i_exotiny.i_rstctl.cnt\[1\] _03136_ net2298 sg13g2_a21oi_1
X_04758_ net1230 _01384_ i_exotiny.i_wb_qspi_mem.cnt_r\[2\] _01509_ VPWR VGND sg13g2_nor3_1
X_04689_ i_exotiny._0315_\[29\] i_exotiny._0314_\[29\] net1271 _01447_ VPWR VGND sg13g2_mux2_1
X_09216_ net763 VGND VPWR _01271_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[6\]
+ clknet_leaf_135_clk_regs sg13g2_dfrbpq_1
X_07477_ _03104_ _01499_ i_exotiny._1266_ VPWR VGND sg13g2_nand2_1
X_08440__245 VPWR VGND net245 sg13g2_tiehi
X_06428_ VPWR _00519_ net3776 VGND sg13g2_inv_1
X_06359_ net2292 net2283 net1031 _00489_ VPWR VGND sg13g2_mux2_1
X_09147_ net835 VGND VPWR _01202_ i_exotiny._0027_\[3\] clknet_leaf_149_clk_regs sg13g2_dfrbpq_2
X_09078_ net1324 VGND VPWR _01133_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[18\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_30_45 VPWR VGND sg13g2_fill_1
X_08029_ net665 VGND VPWR _00110_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[30\]
+ clknet_leaf_61_clk_regs sg13g2_dfrbpq_1
Xhold771 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[10\]
+ VPWR VGND net2598 sg13g2_dlygate4sd3_1
Xhold782 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[8\]
+ VPWR VGND net2609 sg13g2_dlygate4sd3_1
XFILLER_2_936 VPWR VGND sg13g2_decap_8
Xhold760 _00181_ VPWR VGND net2587 sg13g2_dlygate4sd3_1
XFILLER_104_853 VPWR VGND sg13g2_decap_8
Xhold793 _00264_ VPWR VGND net2620 sg13g2_dlygate4sd3_1
XFILLER_77_704 VPWR VGND sg13g2_fill_1
XFILLER_103_374 VPWR VGND sg13g2_decap_8
X_08712__1276 VPWR VGND net1696 sg13g2_tiehi
Xhold1460 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[22\]
+ VPWR VGND net3287 sg13g2_dlygate4sd3_1
Xhold1471 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[14\]
+ VPWR VGND net3298 sg13g2_dlygate4sd3_1
Xhold1482 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[8\]
+ VPWR VGND net3309 sg13g2_dlygate4sd3_1
Xhold1493 i_exotiny._0032_\[0\] VPWR VGND net3320 sg13g2_dlygate4sd3_1
XFILLER_72_453 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_182_clk_regs clknet_5_0__leaf_clk_regs clknet_leaf_182_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_33_818 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_111_clk_regs clknet_5_25__leaf_clk_regs clknet_leaf_111_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_71_63 VPWR VGND sg13g2_fill_2
X_08934__1048 VPWR VGND net1468 sg13g2_tiehi
XFILLER_4_251 VPWR VGND sg13g2_fill_1
XFILLER_99_339 VPWR VGND sg13g2_decap_8
XFILLER_5_796 VPWR VGND sg13g2_decap_4
XFILLER_96_93 VPWR VGND sg13g2_fill_1
X_05730_ _02368_ _02367_ i_exotiny.i_wb_spi.cnt_hbit_r\[4\] VPWR VGND sg13g2_nand2b_1
X_05661_ VGND VPWR i_exotiny._1614_\[3\] net1122 _02317_ _02316_ sg13g2_a21oi_1
X_04612_ VPWR _01374_ _00017_ VGND sg13g2_inv_1
X_08380_ net298 VGND VPWR net2950 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[18\]
+ clknet_leaf_134_clk_regs sg13g2_dfrbpq_1
X_07400_ net1214 VPWR _03052_ VGND _02999_ _03051_ sg13g2_o21ai_1
XFILLER_91_1022 VPWR VGND sg13g2_decap_8
X_05592_ VGND VPWR _02050_ _02265_ _02266_ _02048_ sg13g2_a21oi_1
X_07331_ _02995_ i_exotiny._0369_\[5\] _02994_ VPWR VGND sg13g2_nand2_1
XFILLER_84_0 VPWR VGND sg13g2_fill_2
X_07262_ net2398 net3126 net1006 _00985_ VPWR VGND sg13g2_mux2_1
X_06213_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[25\]
+ net2369 net946 _00368_ VPWR VGND sg13g2_mux2_1
X_07193_ net3589 net3576 net1093 _00929_ VPWR VGND sg13g2_mux2_1
X_09001_ net1401 VGND VPWR _01059_ i_exotiny._1160_\[22\] clknet_leaf_162_clk_regs
+ sg13g2_dfrbpq_1
X_06144_ _02529_ net2682 net1046 _00311_ VPWR VGND sg13g2_mux2_1
X_06075_ net2791 net3091 net956 _00251_ VPWR VGND sg13g2_mux2_1
XFILLER_104_138 VPWR VGND sg13g2_decap_8
X_05026_ net1235 _01756_ _01757_ _01758_ VPWR VGND sg13g2_nor3_2
XFILLER_101_801 VPWR VGND sg13g2_decap_8
XFILLER_99_884 VPWR VGND sg13g2_decap_8
XFILLER_98_383 VPWR VGND sg13g2_decap_8
XFILLER_100_311 VPWR VGND sg13g2_decap_8
XFILLER_58_225 VPWR VGND sg13g2_fill_2
XFILLER_101_878 VPWR VGND sg13g2_decap_8
XFILLER_86_578 VPWR VGND sg13g2_fill_1
XFILLER_74_729 VPWR VGND sg13g2_fill_2
X_06977_ net2280 net2945 net1020 _00750_ VPWR VGND sg13g2_mux2_1
XFILLER_100_388 VPWR VGND sg13g2_decap_8
X_05928_ net2509 _02482_ net973 _00142_ VPWR VGND sg13g2_mux2_1
X_08716_ net1692 VGND VPWR _00774_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[11\]
+ clknet_leaf_117_clk_regs sg13g2_dfrbpq_1
XFILLER_39_494 VPWR VGND sg13g2_fill_2
XFILLER_54_464 VPWR VGND sg13g2_fill_1
X_08647_ net1750 VGND VPWR net3033 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[16\]
+ clknet_leaf_146_clk_regs sg13g2_dfrbpq_1
X_05859_ VGND VPWR _01980_ _02266_ _02447_ _02446_ sg13g2_a21oi_1
XFILLER_82_784 VPWR VGND sg13g2_fill_1
X_08578_ net1826 VGND VPWR net1975 i_exotiny._0314_\[23\] clknet_leaf_180_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_50_670 VPWR VGND sg13g2_fill_1
X_07529_ _03125_ _03106_ _03124_ VPWR VGND sg13g2_nand2b_1
X_08047__647 VPWR VGND net647 sg13g2_tiehi
XFILLER_10_512 VPWR VGND sg13g2_fill_2
XFILLER_104_650 VPWR VGND sg13g2_decap_8
X_08093__601 VPWR VGND net601 sg13g2_tiehi
Xhold590 _00384_ VPWR VGND net2417 sg13g2_dlygate4sd3_1
XFILLER_103_171 VPWR VGND sg13g2_decap_8
XFILLER_66_63 VPWR VGND sg13g2_fill_1
XFILLER_65_729 VPWR VGND sg13g2_fill_2
X_07946__90 VPWR VGND net90 sg13g2_tiehi
Xhold1290 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[31\]
+ VPWR VGND net3117 sg13g2_dlygate4sd3_1
XFILLER_45_486 VPWR VGND sg13g2_decap_4
XFILLER_32_136 VPWR VGND sg13g2_fill_2
X_08423__262 VPWR VGND net262 sg13g2_tiehi
XFILLER_12_1023 VPWR VGND sg13g2_decap_4
X_06900_ VPWR _00695_ _02901_ VGND sg13g2_inv_1
XFILLER_96_865 VPWR VGND sg13g2_decap_8
XFILLER_95_342 VPWR VGND sg13g2_decap_8
X_07880_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[18\]
+ net2259 net982 _01347_ VPWR VGND sg13g2_mux2_1
X_08430__255 VPWR VGND net255 sg13g2_tiehi
X_06831_ net3697 net1096 _02847_ VPWR VGND sg13g2_nor2_1
XFILLER_95_386 VPWR VGND sg13g2_fill_2
X_06762_ _02788_ net1870 net1183 VPWR VGND sg13g2_nand2_1
XFILLER_36_420 VPWR VGND sg13g2_fill_1
X_08501_ net179 VGND VPWR _00575_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[21\]
+ clknet_leaf_71_clk_regs sg13g2_dfrbpq_1
XFILLER_64_762 VPWR VGND sg13g2_fill_2
X_05713_ net1899 net1059 _02356_ VPWR VGND sg13g2_nor2_1
X_08432_ net253 VGND VPWR net2523 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[31\]
+ clknet_leaf_96_clk_regs sg13g2_dfrbpq_1
X_06693_ VPWR VGND _02729_ _02727_ _02728_ i_exotiny.i_wdg_top.o_wb_dat\[0\] _02730_
+ net1181 sg13g2_a221oi_1
XFILLER_36_464 VPWR VGND sg13g2_fill_2
X_05644_ net1124 net1909 _02304_ VPWR VGND sg13g2_nor2b_1
XFILLER_51_467 VPWR VGND sg13g2_fill_1
X_08363_ net315 VGND VPWR net2466 i_exotiny._0014_\[1\] clknet_leaf_140_clk_regs sg13g2_dfrbpq_2
X_05575_ _01385_ _01439_ _02255_ VPWR VGND sg13g2_nor2_1
X_08294_ net384 VGND VPWR net3456 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[28\]
+ clknet_leaf_103_clk_regs sg13g2_dfrbpq_1
X_07314_ net1251 net3768 net1151 _01026_ VPWR VGND sg13g2_mux2_1
X_07245_ net2878 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[8\]
+ net1004 _00968_ VPWR VGND sg13g2_mux2_1
X_07176_ _02951_ net2861 net1011 _00921_ VPWR VGND sg13g2_mux2_1
XFILLER_106_937 VPWR VGND sg13g2_decap_8
XFILLER_105_403 VPWR VGND sg13g2_decap_8
X_06127_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[18\]
+ net3450 net1045 _00296_ VPWR VGND sg13g2_mux2_1
X_06058_ net2271 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[26\]
+ net962 _00243_ VPWR VGND sg13g2_mux2_1
X_05009_ _01701_ _01740_ _01697_ _01741_ VPWR VGND sg13g2_nand3_1
XFILLER_59_523 VPWR VGND sg13g2_fill_1
XFILLER_87_898 VPWR VGND sg13g2_fill_2
XFILLER_86_375 VPWR VGND sg13g2_fill_2
XFILLER_59_589 VPWR VGND sg13g2_fill_1
XFILLER_98_1028 VPWR VGND sg13g2_fill_1
XFILLER_100_196 VPWR VGND sg13g2_decap_8
XFILLER_43_935 VPWR VGND sg13g2_fill_1
XFILLER_11_854 VPWR VGND sg13g2_fill_1
X_08992__990 VPWR VGND net1410 sg13g2_tiehi
XFILLER_7_858 VPWR VGND sg13g2_decap_8
X_08377__301 VPWR VGND net301 sg13g2_tiehi
XFILLER_78_810 VPWR VGND sg13g2_fill_2
X_08866__1120 VPWR VGND net1540 sg13g2_tiehi
X_08884__1098 VPWR VGND net1518 sg13g2_tiehi
XFILLER_92_312 VPWR VGND sg13g2_fill_2
X_09197__784 VPWR VGND net784 sg13g2_tiehi
XFILLER_93_868 VPWR VGND sg13g2_fill_1
XFILLER_92_367 VPWR VGND sg13g2_fill_1
XFILLER_46_740 VPWR VGND sg13g2_fill_2
XFILLER_45_283 VPWR VGND sg13g2_fill_1
XFILLER_60_242 VPWR VGND sg13g2_decap_4
X_05360_ i_exotiny._2034_\[9\] _00023_ _02082_ VPWR VGND sg13g2_xor2_1
X_05291_ _02017_ _01650_ i_exotiny._0016_\[0\] _01641_ i_exotiny._0035_\[0\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_61_2 VPWR VGND sg13g2_fill_1
X_07030_ net3452 net875 _02928_ _02933_ VPWR VGND sg13g2_mux2_1
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_102_406 VPWR VGND sg13g2_decap_8
X_08981_ net1421 VGND VPWR _01039_ i_exotiny._1160_\[2\] clknet_leaf_164_clk_regs
+ sg13g2_dfrbpq_1
X_07932_ net716 VGND VPWR net1921 i_exotiny._1924_\[25\] clknet_leaf_31_clk_regs sg13g2_dfrbpq_1
X_08037__657 VPWR VGND net657 sg13g2_tiehi
X_07863_ i_exotiny._0021_\[1\] net2371 net980 _01330_ VPWR VGND sg13g2_mux2_1
X_06814_ VGND VPWR net1097 _02831_ _00678_ _02832_ sg13g2_a21oi_1
X_07794_ net2071 net2935 net893 _01273_ VPWR VGND sg13g2_mux2_1
X_06745_ VGND VPWR _01411_ net1190 _02774_ net1169 sg13g2_a21oi_1
X_06676_ i_exotiny._0327_\[0\] _01464_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[1\]
+ _02713_ VPWR VGND _01532_ sg13g2_nand4_1
X_08415_ net270 VGND VPWR _00489_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[14\]
+ clknet_leaf_90_clk_regs sg13g2_dfrbpq_1
X_05627_ net1124 net1895 _02291_ VPWR VGND sg13g2_nor2b_1
XFILLER_51_264 VPWR VGND sg13g2_fill_1
X_08083__611 VPWR VGND net611 sg13g2_tiehi
X_08346_ net332 VGND VPWR _00427_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[16\]
+ clknet_leaf_95_clk_regs sg13g2_dfrbpq_1
X_05558_ _02238_ VPWR i_exotiny._1611_\[30\] VGND net1074 _02240_ sg13g2_o21ai_1
X_08277_ net401 VGND VPWR net3480 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[11\]
+ clknet_leaf_100_clk_regs sg13g2_dfrbpq_1
XFILLER_20_662 VPWR VGND sg13g2_fill_1
X_05489_ VGND VPWR i_exotiny._0314_\[2\] net1277 _02187_ _02186_ sg13g2_a21oi_1
X_07228_ net3663 i_exotiny.i_wb_spi.dat_rx_r\[25\] net1086 _00953_ VPWR VGND sg13g2_mux2_1
XFILLER_4_806 VPWR VGND sg13g2_decap_8
XFILLER_106_734 VPWR VGND sg13g2_decap_8
XFILLER_105_200 VPWR VGND sg13g2_decap_8
X_08647__1330 VPWR VGND net1750 sg13g2_tiehi
X_07159_ net3167 net2323 net1011 _00907_ VPWR VGND sg13g2_mux2_1
XFILLER_105_277 VPWR VGND sg13g2_decap_8
Xfanout1106 i_exotiny._2160_ net1106 VPWR VGND sg13g2_buf_1
Xfanout1117 net1120 net1117 VPWR VGND sg13g2_buf_1
Xfanout1128 net1136 net1128 VPWR VGND sg13g2_buf_8
XFILLER_102_951 VPWR VGND sg13g2_decap_8
XFILLER_101_450 VPWR VGND sg13g2_decap_8
X_08090__604 VPWR VGND net604 sg13g2_tiehi
Xfanout1139 net1141 net1139 VPWR VGND sg13g2_buf_8
X_08413__272 VPWR VGND net272 sg13g2_tiehi
XFILLER_86_183 VPWR VGND sg13g2_fill_2
XFILLER_103_60 VPWR VGND sg13g2_fill_2
XFILLER_90_827 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_89_clk_regs clknet_5_31__leaf_clk_regs clknet_leaf_89_clk_regs VPWR VGND
+ sg13g2_buf_8
Xclkbuf_leaf_18_clk_regs clknet_5_7__leaf_clk_regs clknet_leaf_18_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08420__265 VPWR VGND net265 sg13g2_tiehi
XFILLER_98_916 VPWR VGND sg13g2_decap_8
XFILLER_97_415 VPWR VGND sg13g2_decap_8
XFILLER_88_72 VPWR VGND sg13g2_fill_1
XFILLER_3_872 VPWR VGND sg13g2_decap_8
XFILLER_69_139 VPWR VGND sg13g2_fill_1
XFILLER_77_183 VPWR VGND sg13g2_fill_2
XFILLER_19_4 VPWR VGND sg13g2_fill_2
XFILLER_38_537 VPWR VGND sg13g2_fill_1
X_04860_ _01571_ _01576_ _01594_ VPWR VGND sg13g2_and2_1
XFILLER_65_345 VPWR VGND sg13g2_fill_2
XFILLER_38_559 VPWR VGND sg13g2_decap_4
XFILLER_65_389 VPWR VGND sg13g2_fill_2
X_04791_ _01541_ net1283 net1264 VPWR VGND sg13g2_nand2_1
X_06530_ net2224 net2943 net930 _00605_ VPWR VGND sg13g2_mux2_1
X_06461_ net3322 net3342 net937 _00548_ VPWR VGND sg13g2_mux2_1
X_08725__1263 VPWR VGND net1683 sg13g2_tiehi
X_05412_ i_exotiny._2034_\[8\] _02121_ _02123_ VPWR VGND sg13g2_and2_1
X_08200_ net477 VGND VPWR _00281_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[31\]
+ clknet_leaf_69_clk_regs sg13g2_dfrbpq_1
XFILLER_22_949 VPWR VGND sg13g2_fill_1
XFILLER_105_1021 VPWR VGND sg13g2_decap_8
X_09180_ net801 VGND VPWR _01235_ i_exotiny._0026_\[2\] clknet_leaf_79_clk_regs sg13g2_dfrbpq_2
X_06392_ _02574_ _02578_ _02579_ VPWR VGND sg13g2_nor2_1
X_08131_ net1177 VGND VPWR net3560 _00019_ clknet_leaf_36_clk_regs sg13g2_dfrbpq_2
X_05343_ VGND VPWR _01905_ _01907_ _02067_ _01900_ sg13g2_a21oi_1
X_08062_ net632 VGND VPWR net2431 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[31\]
+ clknet_leaf_50_clk_regs sg13g2_dfrbpq_1
X_05274_ _01996_ _01999_ _02000_ VPWR VGND sg13g2_nor2_1
X_08620__1356 VPWR VGND net1776 sg13g2_tiehi
X_07013_ net2075 net2746 net921 _00780_ VPWR VGND sg13g2_mux2_1
XFILLER_102_203 VPWR VGND sg13g2_decap_8
X_08947__1035 VPWR VGND net1455 sg13g2_tiehi
XFILLER_0_319 VPWR VGND sg13g2_fill_1
XFILLER_103_748 VPWR VGND sg13g2_decap_8
X_08964_ net1438 VGND VPWR _01022_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[30\]
+ clknet_leaf_74_clk_regs sg13g2_dfrbpq_1
Xhold1801 _03160_ VPWR VGND net3628 sg13g2_dlygate4sd3_1
X_07915_ net733 VGND VPWR net1942 i_exotiny._1924_\[8\] clknet_leaf_35_clk_regs sg13g2_dfrbpq_1
XFILLER_97_982 VPWR VGND sg13g2_decap_8
Xhold1823 _03178_ VPWR VGND net3650 sg13g2_dlygate4sd3_1
Xhold1812 _00952_ VPWR VGND net3639 sg13g2_dlygate4sd3_1
X_08895_ net1507 VGND VPWR net3664 i_exotiny.i_wb_spi.dat_rx_r\[25\] clknet_leaf_63_clk_regs
+ sg13g2_dfrbpq_1
Xhold1845 i_exotiny._1619_\[2\] VPWR VGND net3672 sg13g2_dlygate4sd3_1
Xhold1834 i_exotiny._0315_\[16\] VPWR VGND net3661 sg13g2_dlygate4sd3_1
Xhold1856 _02913_ VPWR VGND net3683 sg13g2_dlygate4sd3_1
Xhold1878 i_exotiny._1623_ VPWR VGND net3705 sg13g2_dlygate4sd3_1
Xhold1867 i_exotiny._1311_ VPWR VGND net3694 sg13g2_dlygate4sd3_1
X_07846_ net3252 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[22\]
+ net985 _01319_ VPWR VGND sg13g2_mux2_1
X_07777_ _03212_ net3007 net990 _01261_ VPWR VGND sg13g2_mux2_1
Xhold1889 _00073_ VPWR VGND net3716 sg13g2_dlygate4sd3_1
X_08367__311 VPWR VGND net311 sg13g2_tiehi
XFILLER_25_710 VPWR VGND sg13g2_fill_2
X_04989_ _01393_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data[0]
+ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data[0]
+ _01713_ _01718_ _01711_ _01721_ VPWR VGND sg13g2_mux4_1
X_06728_ VPWR VGND net8 _02759_ _02747_ net3795 _02760_ net1182 sg13g2_a221oi_1
XFILLER_25_776 VPWR VGND sg13g2_fill_2
X_06659_ _02698_ _02453_ _02688_ _02699_ VPWR VGND sg13g2_mux2_1
XFILLER_12_448 VPWR VGND sg13g2_fill_2
X_08329_ net349 VGND VPWR net2641 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[31\]
+ clknet_leaf_72_clk_regs sg13g2_dfrbpq_1
X_09276__69 VPWR VGND net69 sg13g2_tiehi
XFILLER_20_481 VPWR VGND sg13g2_fill_2
X_08374__304 VPWR VGND net304 sg13g2_tiehi
XFILLER_4_614 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_136_clk_regs clknet_5_21__leaf_clk_regs clknet_leaf_136_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_106_531 VPWR VGND sg13g2_decap_8
X_09187__794 VPWR VGND net794 sg13g2_tiehi
XFILLER_4_658 VPWR VGND sg13g2_fill_1
XFILLER_4_669 VPWR VGND sg13g2_fill_2
XFILLER_3_146 VPWR VGND sg13g2_fill_1
X_08803__1185 VPWR VGND net1605 sg13g2_tiehi
XFILLER_95_919 VPWR VGND sg13g2_decap_8
XFILLER_0_875 VPWR VGND sg13g2_decap_8
XFILLER_94_429 VPWR VGND sg13g2_fill_1
Xhold8 i_exotiny.i_wb_spi.state_r\[14\] VPWR VGND net1835 sg13g2_dlygate4sd3_1
XFILLER_88_993 VPWR VGND sg13g2_decap_8
XFILLER_16_721 VPWR VGND sg13g2_fill_1
X_09194__787 VPWR VGND net787 sg13g2_tiehi
XFILLER_71_860 VPWR VGND sg13g2_fill_1
XFILLER_43_562 VPWR VGND sg13g2_fill_2
XFILLER_30_212 VPWR VGND sg13g2_fill_1
XFILLER_12_960 VPWR VGND sg13g2_decap_8
XFILLER_30_278 VPWR VGND sg13g2_fill_2
X_08027__667 VPWR VGND net667 sg13g2_tiehi
Xhold408 _00164_ VPWR VGND net2235 sg13g2_dlygate4sd3_1
XFILLER_8_986 VPWR VGND sg13g2_decap_8
Xhold419 _01008_ VPWR VGND net2246 sg13g2_dlygate4sd3_1
X_08073__621 VPWR VGND net621 sg13g2_tiehi
XFILLER_86_908 VPWR VGND sg13g2_fill_1
XFILLER_97_289 VPWR VGND sg13g2_decap_8
X_05961_ net2729 net2477 net966 _00170_ VPWR VGND sg13g2_mux2_1
Xhold1108 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[12\]
+ VPWR VGND net2935 sg13g2_dlygate4sd3_1
X_07700_ net2209 _03198_ net998 _01198_ VPWR VGND sg13g2_mux2_1
Xhold1119 i_exotiny._0013_\[1\] VPWR VGND net2946 sg13g2_dlygate4sd3_1
XFILLER_94_941 VPWR VGND sg13g2_decap_8
X_05892_ _02477_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[4\] VPWR VGND
+ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[3\] sg13g2_nand2b_2
X_08680_ net1728 VGND VPWR net3248 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[7\]
+ clknet_leaf_104_clk_regs sg13g2_dfrbpq_1
X_04912_ _01644_ net1256 _01643_ VPWR VGND sg13g2_nand2_2
X_04843_ _01578_ net1118 _01583_ VPWR VGND sg13g2_and2_1
XFILLER_65_153 VPWR VGND sg13g2_fill_1
X_07631_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[4\]
+ net2097 net899 _01139_ VPWR VGND sg13g2_mux2_1
X_07562_ net3520 net3724 _02178_ _03146_ VPWR VGND sg13g2_nor3_1
X_06513_ i_exotiny._0043_\[2\] net3094 net930 _00588_ VPWR VGND sg13g2_mux2_1
X_09301_ net1535 VGND VPWR _01356_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[27\]
+ clknet_leaf_167_clk_regs sg13g2_dfrbpq_1
X_04774_ _01523_ _01524_ _01525_ VPWR VGND sg13g2_and2_1
X_07493_ VGND VPWR _01386_ net906 _01076_ _03113_ sg13g2_a21oi_1
X_09232_ net747 VGND VPWR _01287_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[22\]
+ clknet_leaf_135_clk_regs sg13g2_dfrbpq_1
X_06444_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[13\]
+ net2232 net934 _00531_ VPWR VGND sg13g2_mux2_1
X_08080__614 VPWR VGND net614 sg13g2_tiehi
X_06375_ i_exotiny._0035_\[1\] net884 _02565_ _02568_ VPWR VGND sg13g2_mux2_1
X_09163_ net819 VGND VPWR _01218_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[19\]
+ clknet_leaf_173_clk_regs sg13g2_dfrbpq_1
X_08403__282 VPWR VGND net282 sg13g2_tiehi
X_05326_ _02041_ VPWR _02050_ VGND _02045_ _02046_ sg13g2_o21ai_1
X_08114_ net580 VGND VPWR _00195_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[19\]
+ clknet_leaf_125_clk_regs sg13g2_dfrbpq_1
X_09094_ net1308 VGND VPWR net3339 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[14\]
+ clknet_leaf_144_clk_regs sg13g2_dfrbpq_1
X_08045_ net649 VGND VPWR net2352 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[14\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
Xhold920 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[25\]
+ VPWR VGND net2747 sg13g2_dlygate4sd3_1
X_05257_ _01983_ _01424_ _01710_ VPWR VGND sg13g2_nand2_1
Xhold931 i_exotiny._0013_\[3\] VPWR VGND net2758 sg13g2_dlygate4sd3_1
Xhold953 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[19\]
+ VPWR VGND net2780 sg13g2_dlygate4sd3_1
Xhold942 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[26\]
+ VPWR VGND net2769 sg13g2_dlygate4sd3_1
Xhold964 i_exotiny._0038_\[1\] VPWR VGND net2791 sg13g2_dlygate4sd3_1
X_05188_ VGND VPWR _01371_ _01739_ _01916_ _01915_ sg13g2_a21oi_1
Xhold986 _00172_ VPWR VGND net2813 sg13g2_dlygate4sd3_1
Xhold975 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[6\]
+ VPWR VGND net2802 sg13g2_dlygate4sd3_1
Xhold997 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[10\]
+ VPWR VGND net2824 sg13g2_dlygate4sd3_1
X_08947_ net1455 VGND VPWR _01005_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[13\]
+ clknet_leaf_54_clk_regs sg13g2_dfrbpq_1
XFILLER_76_418 VPWR VGND sg13g2_fill_2
X_08878_ net1524 VGND VPWR net1969 i_exotiny.i_wb_spi.dat_rx_r\[8\] clknet_leaf_58_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_69_492 VPWR VGND sg13g2_fill_1
Xhold1653 _00358_ VPWR VGND net3480 sg13g2_dlygate4sd3_1
Xhold1620 i_exotiny._0314_\[16\] VPWR VGND net3447 sg13g2_dlygate4sd3_1
Xhold1631 i_exotiny._1611_\[10\] VPWR VGND net3458 sg13g2_dlygate4sd3_1
Xhold1642 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[2\] VPWR
+ VGND net3469 sg13g2_dlygate4sd3_1
X_08410__275 VPWR VGND net275 sg13g2_tiehi
XFILLER_85_985 VPWR VGND sg13g2_decap_8
Xhold1675 _00684_ VPWR VGND net3502 sg13g2_dlygate4sd3_1
XFILLER_56_164 VPWR VGND sg13g2_fill_2
Xhold1686 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[28\]
+ VPWR VGND net3513 sg13g2_dlygate4sd3_1
Xhold1664 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[5\]
+ VPWR VGND net3491 sg13g2_dlygate4sd3_1
X_07829_ net3124 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[5\]
+ net986 _01302_ VPWR VGND sg13g2_mux2_1
XFILLER_72_635 VPWR VGND sg13g2_fill_1
Xhold1697 i_exotiny._1489_\[0\] VPWR VGND net3524 sg13g2_dlygate4sd3_1
XFILLER_40_521 VPWR VGND sg13g2_decap_4
XFILLER_13_768 VPWR VGND sg13g2_fill_2
XFILLER_44_99 VPWR VGND sg13g2_decap_8
XFILLER_9_739 VPWR VGND sg13g2_fill_1
XFILLER_5_945 VPWR VGND sg13g2_decap_8
XFILLER_4_411 VPWR VGND sg13g2_fill_2
XFILLER_4_455 VPWR VGND sg13g2_fill_1
XFILLER_48_654 VPWR VGND sg13g2_fill_1
XFILLER_48_632 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_33_clk_regs clknet_5_8__leaf_clk_regs clknet_leaf_33_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_78_1026 VPWR VGND sg13g2_fill_2
XFILLER_91_966 VPWR VGND sg13g2_decap_8
XFILLER_93_5 VPWR VGND sg13g2_fill_2
X_06160_ net3191 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[12\]
+ net953 _00322_ VPWR VGND sg13g2_mux2_1
Xhold216 _00211_ VPWR VGND net2043 sg13g2_dlygate4sd3_1
Xhold205 _00042_ VPWR VGND net2032 sg13g2_dlygate4sd3_1
X_08357__321 VPWR VGND net321 sg13g2_tiehi
X_06091_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[17\]
+ net3279 net955 _00267_ VPWR VGND sg13g2_mux2_1
X_05111_ VGND VPWR _01371_ _01739_ _01841_ _01840_ sg13g2_a21oi_1
Xhold227 i_exotiny.i_wdg_top.clk_div_inst.cnt\[17\] VPWR VGND net2054 sg13g2_dlygate4sd3_1
Xhold238 i_exotiny._1160_\[9\] VPWR VGND net2065 sg13g2_dlygate4sd3_1
Xhold249 _00776_ VPWR VGND net2076 sg13g2_dlygate4sd3_1
X_05042_ net1236 _01753_ _01754_ _01774_ VPWR VGND sg13g2_nor3_2
X_07995__136 VPWR VGND net136 sg13g2_tiehi
X_08801_ net1607 VGND VPWR net3635 i_exotiny.i_wb_spi.state_r\[0\] clknet_leaf_32_clk_regs
+ sg13g2_dfrbpq_2
X_06993_ net2178 _02927_ net1019 _00762_ VPWR VGND sg13g2_mux2_1
X_05944_ net2418 net3460 net969 _00153_ VPWR VGND sg13g2_mux2_1
X_08732_ net1676 VGND VPWR _00790_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[27\]
+ clknet_leaf_118_clk_regs sg13g2_dfrbpq_1
X_08663_ net1203 VGND VPWR i_exotiny._2043_\[0\] i_exotiny._2034_\[0\] net1228 sg13g2_dfrbpq_2
XFILLER_38_142 VPWR VGND sg13g2_fill_2
XFILLER_39_665 VPWR VGND sg13g2_decap_4
XFILLER_39_687 VPWR VGND sg13g2_fill_2
X_05875_ _02462_ _02457_ _02461_ net1184 _01419_ VPWR VGND sg13g2_a22oi_1
X_07614_ _03180_ net3842 net1880 _03176_ VPWR VGND sg13g2_and3_1
X_04826_ net1846 net1858 net1853 net1837 _01566_ VPWR VGND sg13g2_nor4_1
X_08594_ net1802 VGND VPWR _00666_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data[0]
+ clknet_leaf_26_clk_regs sg13g2_dfrbpq_2
X_08897__1085 VPWR VGND net1505 sg13g2_tiehi
X_08364__314 VPWR VGND net314 sg13g2_tiehi
XFILLER_42_819 VPWR VGND sg13g2_fill_2
X_07545_ _03133_ _03135_ _01106_ VPWR VGND sg13g2_nor2_1
X_04757_ net1196 _01446_ net3695 _00005_ VPWR VGND sg13g2_nor3_1
XFILLER_22_543 VPWR VGND sg13g2_fill_1
X_07476_ net1211 net3580 _03021_ _01069_ VPWR VGND sg13g2_a21o_1
X_04688_ i_exotiny._1489_\[3\] i_exotiny._1489_\[0\] _01446_ VPWR VGND sg13g2_and2_1
X_09215_ net764 VGND VPWR _01270_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[5\]
+ clknet_leaf_129_clk_regs sg13g2_dfrbpq_1
X_06427_ net1284 VPWR _02605_ VGND net3775 _02604_ sg13g2_o21ai_1
X_06358_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[17\]
+ net3354 net1028 _00488_ VPWR VGND sg13g2_mux2_1
X_09146_ net836 VGND VPWR _01201_ i_exotiny._0027_\[2\] clknet_leaf_149_clk_regs sg13g2_dfrbpq_2
X_09077_ net1325 VGND VPWR net2056 i_exotiny.i_wdg_top.clk_div_inst.cnt\[17\] clknet_leaf_50_clk_regs
+ sg13g2_dfrbpq_1
X_06289_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[25\]
+ net2367 net940 _00432_ VPWR VGND sg13g2_mux2_1
X_05309_ _02019_ _02024_ _02034_ _02035_ VPWR VGND sg13g2_nor3_2
X_08028_ net666 VGND VPWR net3371 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[29\]
+ clknet_leaf_67_clk_regs sg13g2_dfrbpq_1
XFILLER_2_915 VPWR VGND sg13g2_decap_8
XFILLER_104_832 VPWR VGND sg13g2_decap_8
Xhold750 _00504_ VPWR VGND net2577 sg13g2_dlygate4sd3_1
Xhold772 _00090_ VPWR VGND net2599 sg13g2_dlygate4sd3_1
X_08371__307 VPWR VGND net307 sg13g2_tiehi
Xhold761 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[28\]
+ VPWR VGND net2588 sg13g2_dlygate4sd3_1
X_09184__797 VPWR VGND net797 sg13g2_tiehi
Xhold794 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[16\]
+ VPWR VGND net2621 sg13g2_dlygate4sd3_1
Xhold783 _00530_ VPWR VGND net2610 sg13g2_dlygate4sd3_1
XFILLER_39_11 VPWR VGND sg13g2_decap_8
XFILLER_103_353 VPWR VGND sg13g2_decap_8
X_08684__1304 VPWR VGND net1724 sg13g2_tiehi
Xclkbuf_4_1_0_clk_regs clknet_0_clk_regs clknet_4_1_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_39_99 VPWR VGND sg13g2_decap_4
Xhold1450 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[9\]
+ VPWR VGND net3277 sg13g2_dlygate4sd3_1
Xhold1461 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[15\]
+ VPWR VGND net3288 sg13g2_dlygate4sd3_1
XFILLER_29_131 VPWR VGND sg13g2_fill_2
Xhold1494 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[30\]
+ VPWR VGND net3321 sg13g2_dlygate4sd3_1
X_08017__677 VPWR VGND net677 sg13g2_tiehi
XFILLER_72_421 VPWR VGND sg13g2_fill_1
XFILLER_55_21 VPWR VGND sg13g2_fill_2
Xhold1483 _00735_ VPWR VGND net3310 sg13g2_dlygate4sd3_1
Xhold1472 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[18\]
+ VPWR VGND net3299 sg13g2_dlygate4sd3_1
XFILLER_17_315 VPWR VGND sg13g2_fill_1
XFILLER_45_635 VPWR VGND sg13g2_fill_1
XFILLER_45_646 VPWR VGND sg13g2_decap_4
XFILLER_73_988 VPWR VGND sg13g2_fill_1
XFILLER_60_627 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_151_clk_regs clknet_5_18__leaf_clk_regs clknet_leaf_151_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08063__631 VPWR VGND net631 sg13g2_tiehi
X_08942__1040 VPWR VGND net1460 sg13g2_tiehi
X_09091__891 VPWR VGND net1311 sg13g2_tiehi
XFILLER_99_318 VPWR VGND sg13g2_decap_8
XFILLER_68_705 VPWR VGND sg13g2_fill_2
XFILLER_96_83 VPWR VGND sg13g2_fill_1
XFILLER_95_546 VPWR VGND sg13g2_fill_1
XFILLER_1_992 VPWR VGND sg13g2_decap_8
X_08070__624 VPWR VGND net624 sg13g2_tiehi
XFILLER_36_635 VPWR VGND sg13g2_decap_8
X_05660_ net1122 net1963 _02316_ VPWR VGND sg13g2_nor2b_1
XFILLER_91_1001 VPWR VGND sg13g2_decap_8
X_04611_ VPWR _01373_ _00018_ VGND sg13g2_inv_1
X_05591_ VGND VPWR i_exotiny._0352_ _01831_ _02265_ _02264_ sg13g2_a21oi_1
XFILLER_51_649 VPWR VGND sg13g2_decap_8
XFILLER_50_148 VPWR VGND sg13g2_fill_2
XFILLER_32_841 VPWR VGND sg13g2_fill_1
X_07330_ i_exotiny._0369_\[4\] i_exotiny._0369_\[2\] _02994_ VPWR VGND sg13g2_nor2_1
X_07261_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[28\]
+ net2759 net1003 _00984_ VPWR VGND sg13g2_mux2_1
X_09000_ net1402 VGND VPWR net3536 i_exotiny._1160_\[21\] clknet_leaf_161_clk_regs
+ sg13g2_dfrbpq_1
X_06212_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[24\]
+ net2375 net947 _00367_ VPWR VGND sg13g2_mux2_1
X_07192_ net9 net3589 net1093 _00928_ VPWR VGND sg13g2_mux2_1
X_08762__1226 VPWR VGND net1646 sg13g2_tiehi
X_06143_ i_exotiny._0037_\[1\] net882 _02526_ _02529_ VPWR VGND sg13g2_mux2_1
X_08588__1388 VPWR VGND net1808 sg13g2_tiehi
X_08400__285 VPWR VGND net285 sg13g2_tiehi
XFILLER_105_629 VPWR VGND sg13g2_decap_8
XFILLER_104_117 VPWR VGND sg13g2_decap_8
XFILLER_104_106 VPWR VGND sg13g2_fill_2
X_06074_ net2933 net3461 net957 _00250_ VPWR VGND sg13g2_mux2_1
XFILLER_99_863 VPWR VGND sg13g2_decap_8
X_05025_ _01757_ i_exotiny._0079_\[2\] VPWR VGND i_exotiny._0079_\[3\] sg13g2_nand2b_2
XFILLER_98_362 VPWR VGND sg13g2_decap_8
XFILLER_101_857 VPWR VGND sg13g2_decap_8
XFILLER_59_749 VPWR VGND sg13g2_fill_2
XFILLER_100_367 VPWR VGND sg13g2_decap_8
X_06976_ net2329 net2819 net1022 _00749_ VPWR VGND sg13g2_mux2_1
X_05927_ net876 i_exotiny._0019_\[2\] _02478_ _02482_ VPWR VGND sg13g2_mux2_1
X_08715_ net1693 VGND VPWR net3035 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[10\]
+ clknet_leaf_120_clk_regs sg13g2_dfrbpq_1
XFILLER_82_741 VPWR VGND sg13g2_fill_1
X_08646_ net1751 VGND VPWR net3042 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[15\]
+ clknet_leaf_145_clk_regs sg13g2_dfrbpq_1
X_05858_ _02429_ VPWR _02446_ VGND _01980_ _02266_ sg13g2_o21ai_1
X_04809_ _01485_ _01521_ _01553_ VPWR VGND sg13g2_nor2_2
X_05789_ _02410_ i_exotiny.i_wdg_top.o_wb_dat\[10\] net1144 VPWR VGND sg13g2_nand2_1
X_08577_ net49 VGND VPWR net1966 i_exotiny._0314_\[22\] clknet_leaf_180_clk_regs sg13g2_dfrbpq_1
X_07528_ VPWR VGND _01814_ _01500_ _01752_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[3\]
+ _03124_ _01686_ sg13g2_a221oi_1
X_07459_ VGND VPWR net3637 net1080 _03096_ _03077_ sg13g2_a21oi_1
X_08738__1250 VPWR VGND net1670 sg13g2_tiehi
XFILLER_10_579 VPWR VGND sg13g2_fill_2
X_09129_ net853 VGND VPWR net2195 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[17\]
+ clknet_leaf_154_clk_regs sg13g2_dfrbpq_1
X_09249__558 VPWR VGND net558 sg13g2_tiehi
Xhold580 _00162_ VPWR VGND net2407 sg13g2_dlygate4sd3_1
XFILLER_1_211 VPWR VGND sg13g2_fill_1
XFILLER_2_734 VPWR VGND sg13g2_decap_4
XFILLER_103_150 VPWR VGND sg13g2_decap_8
Xhold591 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[9\]
+ VPWR VGND net2418 sg13g2_dlygate4sd3_1
XFILLER_2_789 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_66_53 VPWR VGND sg13g2_fill_2
XFILLER_65_708 VPWR VGND sg13g2_fill_2
XFILLER_92_549 VPWR VGND sg13g2_fill_1
Xhold1291 _00585_ VPWR VGND net3118 sg13g2_dlygate4sd3_1
Xhold1280 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[15\]
+ VPWR VGND net3107 sg13g2_dlygate4sd3_1
X_08347__331 VPWR VGND net331 sg13g2_tiehi
XFILLER_33_605 VPWR VGND sg13g2_fill_1
XFILLER_9_355 VPWR VGND sg13g2_fill_1
XFILLER_12_1002 VPWR VGND sg13g2_decap_8
X_08354__324 VPWR VGND net324 sg13g2_tiehi
X_08584__1394 VPWR VGND net1814 sg13g2_tiehi
XFILLER_96_844 VPWR VGND sg13g2_decap_8
XFILLER_95_321 VPWR VGND sg13g2_decap_8
XFILLER_95_376 VPWR VGND sg13g2_fill_2
X_06830_ VGND VPWR net3572 net1131 _02846_ _02845_ sg13g2_a21oi_1
X_06761_ VGND VPWR _01506_ _02785_ _00670_ _02787_ sg13g2_a21oi_1
X_08500_ net180 VGND VPWR net2229 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[20\]
+ clknet_leaf_108_clk_regs sg13g2_dfrbpq_1
XFILLER_64_741 VPWR VGND sg13g2_fill_1
XFILLER_64_730 VPWR VGND sg13g2_fill_1
X_05712_ VGND VPWR i_exotiny._1618_\[0\] net1114 _02355_ _02354_ sg13g2_a21oi_1
X_06692_ VGND VPWR _01407_ net1193 _02729_ net1169 sg13g2_a21oi_1
X_08816__1172 VPWR VGND net1592 sg13g2_tiehi
X_05643_ net1922 net1066 _02303_ VPWR VGND sg13g2_nor2_1
X_08431_ net254 VGND VPWR _00505_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[30\]
+ clknet_leaf_96_clk_regs sg13g2_dfrbpq_1
XFILLER_63_284 VPWR VGND sg13g2_fill_1
X_08361__317 VPWR VGND net317 sg13g2_tiehi
X_08362_ net316 VGND VPWR _00443_ i_exotiny._0014_\[0\] clknet_leaf_140_clk_regs sg13g2_dfrbpq_2
X_05574_ net1984 VPWR _02254_ VGND i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[0\]
+ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[1\] sg13g2_o21ai_1
X_08293_ net385 VGND VPWR _00374_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[27\]
+ clknet_leaf_100_clk_regs sg13g2_dfrbpq_1
XFILLER_20_833 VPWR VGND sg13g2_fill_1
X_07313_ net3690 i_exotiny._0369_\[3\] net1150 _01025_ VPWR VGND sg13g2_mux2_1
X_07244_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[11\]
+ net2467 net1006 _00967_ VPWR VGND sg13g2_mux2_1
XFILLER_106_916 VPWR VGND sg13g2_decap_8
X_07175_ net3397 net876 _02947_ _02951_ VPWR VGND sg13g2_mux2_1
X_06126_ net3038 net2979 net1046 _00295_ VPWR VGND sg13g2_mux2_1
XFILLER_105_459 VPWR VGND sg13g2_decap_8
X_06057_ net2795 net3389 net961 _00242_ VPWR VGND sg13g2_mux2_1
X_05008_ _01694_ _01698_ _01689_ _01740_ VPWR VGND sg13g2_nand3_1
XFILLER_98_192 VPWR VGND sg13g2_fill_1
XFILLER_98_1007 VPWR VGND sg13g2_decap_8
XFILLER_47_719 VPWR VGND sg13g2_fill_1
XFILLER_47_708 VPWR VGND sg13g2_decap_8
X_08053__641 VPWR VGND net641 sg13g2_tiehi
X_06959_ i_exotiny._0034_\[1\] net2677 net1018 _00732_ VPWR VGND sg13g2_mux2_1
XFILLER_28_933 VPWR VGND sg13g2_fill_2
XFILLER_46_218 VPWR VGND sg13g2_fill_2
XFILLER_55_752 VPWR VGND sg13g2_fill_2
XFILLER_54_295 VPWR VGND sg13g2_fill_2
X_08629_ net774 VGND VPWR net1986 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[2\]
+ clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
XFILLER_23_671 VPWR VGND sg13g2_fill_1
XFILLER_7_848 VPWR VGND sg13g2_decap_4
X_08060__634 VPWR VGND net634 sg13g2_tiehi
X_09288__1403 VPWR VGND net1823 sg13g2_tiehi
XFILLER_81_1022 VPWR VGND sg13g2_decap_8
X_08569__66 VPWR VGND net66 sg13g2_tiehi
XFILLER_105_993 VPWR VGND sg13g2_decap_8
XFILLER_104_481 VPWR VGND sg13g2_decap_8
XFILLER_96_129 VPWR VGND sg13g2_fill_1
X_08892__1090 VPWR VGND net1510 sg13g2_tiehi
XFILLER_28_9 VPWR VGND sg13g2_fill_1
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_92_324 VPWR VGND sg13g2_fill_2
XFILLER_18_410 VPWR VGND sg13g2_fill_1
Xfanout890 _02444_ net890 VPWR VGND sg13g2_buf_8
XFILLER_92_357 VPWR VGND sg13g2_fill_1
XFILLER_19_999 VPWR VGND sg13g2_fill_2
XFILLER_60_298 VPWR VGND sg13g2_fill_1
X_05290_ _02016_ _01638_ i_exotiny._0029_\[0\] _01626_ i_exotiny._0014_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_08497__183 VPWR VGND net183 sg13g2_tiehi
X_08980_ net1422 VGND VPWR net2045 i_exotiny._1160_\[1\] clknet_leaf_18_clk_regs sg13g2_dfrbpq_1
XFILLER_68_321 VPWR VGND sg13g2_fill_2
X_07931_ net717 VGND VPWR net2529 i_exotiny._1924_\[24\] clknet_leaf_34_clk_regs sg13g2_dfrbpq_1
XFILLER_56_505 VPWR VGND sg13g2_fill_1
X_07862_ i_exotiny._0021_\[0\] net2069 net982 _01329_ VPWR VGND sg13g2_mux2_1
XFILLER_83_324 VPWR VGND sg13g2_fill_1
X_06813_ net3630 net1097 _02832_ VPWR VGND sg13g2_nor2_1
XFILLER_84_858 VPWR VGND sg13g2_fill_2
X_07793_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[7\]
+ net3292 net891 _01272_ VPWR VGND sg13g2_mux2_1
X_06744_ _02773_ net3708 net1183 VPWR VGND sg13g2_nand2_1
XFILLER_37_774 VPWR VGND sg13g2_fill_2
XFILLER_52_733 VPWR VGND sg13g2_fill_2
X_06675_ net1224 net1234 net1249 _02712_ VPWR VGND _01463_ sg13g2_nand4_1
X_08414_ net271 VGND VPWR net3355 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[13\]
+ clknet_leaf_90_clk_regs sg13g2_dfrbpq_1
X_05626_ VGND VPWR net1066 _02290_ _00032_ _02288_ sg13g2_a21oi_1
XFILLER_40_928 VPWR VGND sg13g2_fill_1
X_08345_ net333 VGND VPWR net3406 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[15\]
+ clknet_leaf_98_clk_regs sg13g2_dfrbpq_1
X_05557_ VGND VPWR net3610 net1277 _02240_ _02239_ sg13g2_a21oi_1
X_08276_ net402 VGND VPWR net2428 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[10\]
+ clknet_leaf_102_clk_regs sg13g2_dfrbpq_1
X_05488_ net1279 net1233 _02186_ VPWR VGND sg13g2_nor2b_1
X_07227_ net3638 i_exotiny.i_wb_spi.dat_rx_r\[24\] net1087 _00952_ VPWR VGND sg13g2_mux2_1
XFILLER_106_713 VPWR VGND sg13g2_decap_8
X_07158_ net3016 net3107 net1008 _00906_ VPWR VGND sg13g2_mux2_1
X_06109_ net3169 _02524_ net959 _00281_ VPWR VGND sg13g2_mux2_1
XFILLER_105_256 VPWR VGND sg13g2_decap_8
X_08337__341 VPWR VGND net341 sg13g2_tiehi
XFILLER_65_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
X_07089_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[17\]
+ net2158 net915 _00844_ VPWR VGND sg13g2_mux2_1
XFILLER_102_930 VPWR VGND sg13g2_decap_8
Xfanout1118 net1119 net1118 VPWR VGND sg13g2_buf_8
Xfanout1129 net1136 net1129 VPWR VGND sg13g2_buf_1
Xfanout1107 net1108 net1107 VPWR VGND sg13g2_buf_2
XFILLER_59_343 VPWR VGND sg13g2_fill_1
XFILLER_87_674 VPWR VGND sg13g2_fill_1
X_08869__1114 VPWR VGND net1534 sg13g2_tiehi
XFILLER_70_541 VPWR VGND sg13g2_fill_2
X_08344__334 VPWR VGND net334 sg13g2_tiehi
Xclkbuf_leaf_58_clk_regs clknet_5_14__leaf_clk_regs clknet_leaf_58_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08790__1198 VPWR VGND net1618 sg13g2_tiehi
XFILLER_12_91 VPWR VGND sg13g2_fill_1
XFILLER_3_851 VPWR VGND sg13g2_decap_8
XFILLER_105_790 VPWR VGND sg13g2_decap_8
X_08351__327 VPWR VGND net327 sg13g2_tiehi
XFILLER_69_129 VPWR VGND sg13g2_fill_1
XFILLER_78_696 VPWR VGND sg13g2_fill_2
XFILLER_93_677 VPWR VGND sg13g2_fill_1
XFILLER_53_519 VPWR VGND sg13g2_fill_1
X_04790_ _01538_ _01539_ net1231 _01540_ VPWR VGND sg13g2_nand3_1
XFILLER_46_560 VPWR VGND sg13g2_decap_8
XFILLER_34_722 VPWR VGND sg13g2_fill_1
Xclkbuf_4_14_0_clk_regs clknet_0_clk_regs clknet_4_14_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_22_917 VPWR VGND sg13g2_fill_1
X_06460_ net2249 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[25\]
+ net934 _00547_ VPWR VGND sg13g2_mux2_1
X_05411_ i_exotiny._2034_\[8\] _02121_ _02122_ VPWR VGND sg13g2_nor2_1
XFILLER_105_1000 VPWR VGND sg13g2_decap_8
X_08130_ net1178 VGND VPWR net2043 _00018_ clknet_leaf_35_clk_regs sg13g2_dfrbpq_2
X_06391_ _02577_ VPWR _02578_ VGND net1273 _01391_ sg13g2_o21ai_1
X_05342_ _02066_ _01388_ _01818_ VPWR VGND sg13g2_nand2_1
X_08061_ net633 VGND VPWR net2510 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[30\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
XFILLER_88_1028 VPWR VGND sg13g2_fill_1
X_05273_ _01992_ _01997_ _01990_ _01999_ VPWR VGND _01998_ sg13g2_nand4_1
X_08043__651 VPWR VGND net651 sg13g2_tiehi
X_07012_ net2645 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[20\]
+ net922 _00779_ VPWR VGND sg13g2_mux2_1
XFILLER_103_705 VPWR VGND sg13g2_fill_2
XFILLER_103_727 VPWR VGND sg13g2_decap_8
X_08963_ net1439 VGND VPWR _01021_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[29\]
+ clknet_leaf_61_clk_regs sg13g2_dfrbpq_1
XFILLER_102_259 VPWR VGND sg13g2_decap_8
XFILLER_97_961 VPWR VGND sg13g2_decap_8
Xhold1802 _01119_ VPWR VGND net3629 sg13g2_dlygate4sd3_1
X_07914_ net734 VGND VPWR net1896 i_exotiny._1924_\[7\] clknet_leaf_34_clk_regs sg13g2_dfrbpq_1
Xhold1813 i_exotiny.i_wb_spi.state_r\[0\] VPWR VGND net3640 sg13g2_dlygate4sd3_1
X_08894_ net1508 VGND VPWR net3639 i_exotiny.i_wb_spi.dat_rx_r\[24\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_1
Xhold1824 i_exotiny._1793_ VPWR VGND net3651 sg13g2_dlygate4sd3_1
Xhold1835 _01086_ VPWR VGND net3662 sg13g2_dlygate4sd3_1
Xhold1846 _00690_ VPWR VGND net3673 sg13g2_dlygate4sd3_1
Xhold1868 _01508_ VPWR VGND net3695 sg13g2_dlygate4sd3_1
X_07845_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[25\]
+ net2347 net985 _01318_ VPWR VGND sg13g2_mux2_1
Xhold1857 i_exotiny._0590_ VPWR VGND net3684 sg13g2_dlygate4sd3_1
X_08050__644 VPWR VGND net644 sg13g2_tiehi
X_07776_ i_exotiny._0026_\[0\] net888 _03210_ _03212_ VPWR VGND sg13g2_mux2_1
Xhold1879 i_exotiny._0315_\[17\] VPWR VGND net3706 sg13g2_dlygate4sd3_1
X_04988_ VGND VPWR _01365_ _01712_ _01720_ _01719_ sg13g2_a21oi_1
X_06727_ VGND VPWR _01408_ net1193 _02759_ _02758_ sg13g2_a21oi_1
X_08857__1129 VPWR VGND net1549 sg13g2_tiehi
X_06658_ _02698_ _02259_ _02697_ VPWR VGND sg13g2_nand2_1
X_05609_ net1903 net1067 _02278_ VPWR VGND sg13g2_nor2_1
X_06589_ net3382 net1162 _02649_ VPWR VGND sg13g2_nor2_1
X_08328_ net350 VGND VPWR _00409_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[30\]
+ clknet_leaf_73_clk_regs sg13g2_dfrbpq_1
X_08259_ net418 VGND VPWR _00340_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[26\]
+ clknet_leaf_49_clk_regs sg13g2_dfrbpq_1
XFILLER_106_510 VPWR VGND sg13g2_decap_8
XFILLER_106_587 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_176_clk_regs clknet_5_1__leaf_clk_regs clknet_leaf_176_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_88_972 VPWR VGND sg13g2_decap_8
XFILLER_58_54 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_105_clk_regs clknet_5_22__leaf_clk_regs clknet_leaf_105_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_0_854 VPWR VGND sg13g2_decap_8
X_08775__1213 VPWR VGND net1633 sg13g2_tiehi
Xhold9 _00873_ VPWR VGND net1836 sg13g2_dlygate4sd3_1
XFILLER_58_76 VPWR VGND sg13g2_fill_2
XFILLER_75_644 VPWR VGND sg13g2_fill_1
X_08487__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_31_769 VPWR VGND sg13g2_fill_1
XFILLER_8_965 VPWR VGND sg13g2_decap_8
Xhold409 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[24\]
+ VPWR VGND net2236 sg13g2_dlygate4sd3_1
XFILLER_99_83 VPWR VGND sg13g2_fill_1
X_08494__186 VPWR VGND net186 sg13g2_tiehi
XFILLER_97_268 VPWR VGND sg13g2_decap_8
XFILLER_94_920 VPWR VGND sg13g2_decap_8
X_05960_ net2458 net2772 net968 _00169_ VPWR VGND sg13g2_mux2_1
Xhold1109 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[29\]
+ VPWR VGND net2936 sg13g2_dlygate4sd3_1
X_05891_ net1262 _02475_ _02476_ VPWR VGND sg13g2_nor2b_2
X_04911_ _01617_ _01640_ _01643_ VPWR VGND sg13g2_nor2_2
XFILLER_94_997 VPWR VGND sg13g2_decap_8
X_04842_ _01379_ _01570_ _01582_ VPWR VGND sg13g2_and2_1
X_07630_ i_exotiny._0024_\[3\] net2917 net896 _01138_ VPWR VGND sg13g2_mux2_1
X_07561_ net1225 net1231 _03145_ _01112_ VPWR VGND sg13g2_nor3_1
X_08638__1339 VPWR VGND net1759 sg13g2_tiehi
X_04773_ _01524_ net1146 _01513_ VPWR VGND sg13g2_nand2_1
X_06512_ i_exotiny._0043_\[1\] net2285 net932 _00587_ VPWR VGND sg13g2_mux2_1
X_09300_ net1537 VGND VPWR _01355_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[26\]
+ clknet_leaf_171_clk_regs sg13g2_dfrbpq_1
X_08327__351 VPWR VGND net351 sg13g2_tiehi
XFILLER_55_1027 VPWR VGND sg13g2_fill_2
X_07492_ net3537 net906 _03113_ VPWR VGND sg13g2_nor2_1
X_06443_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[12\]
+ net2609 net937 _00530_ VPWR VGND sg13g2_mux2_1
X_09231_ net748 VGND VPWR _01286_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[21\]
+ clknet_leaf_129_clk_regs sg13g2_dfrbpq_1
X_06374_ _02567_ net3324 net1029 _00503_ VPWR VGND sg13g2_mux2_1
X_09162_ net820 VGND VPWR _01217_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[18\]
+ clknet_leaf_148_clk_regs sg13g2_dfrbpq_1
X_08113_ net581 VGND VPWR _00194_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[18\]
+ clknet_leaf_122_clk_regs sg13g2_dfrbpq_1
X_05325_ _02041_ _02045_ _02046_ _02049_ VPWR VGND sg13g2_or3_1
X_09093_ net1309 VGND VPWR _01148_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[13\]
+ clknet_leaf_142_clk_regs sg13g2_dfrbpq_1
X_08044_ net650 VGND VPWR net2884 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[13\]
+ clknet_leaf_54_clk_regs sg13g2_dfrbpq_1
Xhold910 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[16\]
+ VPWR VGND net2737 sg13g2_dlygate4sd3_1
Xhold921 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[21\]
+ VPWR VGND net2748 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_3_clk_regs clknet_5_2__leaf_clk_regs clknet_leaf_3_clk_regs VPWR VGND
+ sg13g2_buf_8
X_05256_ VGND VPWR _01743_ _01981_ _01982_ _01702_ sg13g2_a21oi_1
Xhold943 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[26\]
+ VPWR VGND net2770 sg13g2_dlygate4sd3_1
Xhold932 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[24\]
+ VPWR VGND net2759 sg13g2_dlygate4sd3_1
Xhold954 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[27\]
+ VPWR VGND net2781 sg13g2_dlygate4sd3_1
X_05187_ _01708_ VPWR _01915_ VGND i_exotiny._0315_\[4\] _01424_ sg13g2_o21ai_1
XFILLER_103_535 VPWR VGND sg13g2_decap_8
Xhold965 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[12\]
+ VPWR VGND net2792 sg13g2_dlygate4sd3_1
Xhold987 i_exotiny._0016_\[3\] VPWR VGND net2814 sg13g2_dlygate4sd3_1
Xhold976 i_exotiny._0034_\[2\] VPWR VGND net2803 sg13g2_dlygate4sd3_1
Xhold998 _00592_ VPWR VGND net2825 sg13g2_dlygate4sd3_1
X_08334__344 VPWR VGND net344 sg13g2_tiehi
X_08946_ net1456 VGND VPWR net2716 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[12\]
+ clknet_leaf_75_clk_regs sg13g2_dfrbpq_1
Xhold1610 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[31\]
+ VPWR VGND net3437 sg13g2_dlygate4sd3_1
X_08877_ net1525 VGND VPWR net1936 i_exotiny.i_wb_spi.dat_rx_r\[7\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_1
Xhold1632 i_exotiny._0027_\[3\] VPWR VGND net3459 sg13g2_dlygate4sd3_1
Xhold1621 _00640_ VPWR VGND net3448 sg13g2_dlygate4sd3_1
XFILLER_28_35 VPWR VGND sg13g2_fill_2
Xhold1643 _01499_ VPWR VGND net3470 sg13g2_dlygate4sd3_1
XFILLER_84_441 VPWR VGND sg13g2_fill_2
XFILLER_57_677 VPWR VGND sg13g2_fill_2
Xhold1687 _00204_ VPWR VGND net3514 sg13g2_dlygate4sd3_1
Xhold1676 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[23\]
+ VPWR VGND net3503 sg13g2_dlygate4sd3_1
Xhold1654 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[6\]
+ VPWR VGND net3481 sg13g2_dlygate4sd3_1
Xhold1665 _01298_ VPWR VGND net3492 sg13g2_dlygate4sd3_1
X_07828_ net3119 net2134 net987 _01301_ VPWR VGND sg13g2_mux2_1
XFILLER_56_198 VPWR VGND sg13g2_fill_2
Xhold1698 i_exotiny._0023_\[2\] VPWR VGND net3525 sg13g2_dlygate4sd3_1
X_07759_ net2743 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[11\]
+ net990 _01244_ VPWR VGND sg13g2_mux2_1
XFILLER_53_861 VPWR VGND sg13g2_fill_2
X_08341__337 VPWR VGND net337 sg13g2_tiehi
XFILLER_40_588 VPWR VGND sg13g2_fill_2
XFILLER_5_924 VPWR VGND sg13g2_decap_8
XFILLER_106_384 VPWR VGND sg13g2_decap_8
XFILLER_76_986 VPWR VGND sg13g2_fill_1
XFILLER_36_817 VPWR VGND sg13g2_fill_1
XFILLER_91_945 VPWR VGND sg13g2_decap_8
X_08033__661 VPWR VGND net661 sg13g2_tiehi
XFILLER_47_176 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_73_clk_regs clknet_5_24__leaf_clk_regs clknet_leaf_73_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_62_135 VPWR VGND sg13g2_fill_2
XFILLER_90_477 VPWR VGND sg13g2_fill_2
XFILLER_44_883 VPWR VGND sg13g2_fill_1
XFILLER_43_382 VPWR VGND sg13g2_fill_2
XFILLER_86_5 VPWR VGND sg13g2_fill_1
XFILLER_8_740 VPWR VGND sg13g2_fill_1
XFILLER_102_1014 VPWR VGND sg13g2_decap_8
X_05110_ _01708_ VPWR _01840_ VGND i_exotiny._0315_\[4\] _01425_ sg13g2_o21ai_1
Xhold206 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.genblk7.g_value.r_value[0]
+ VPWR VGND net2033 sg13g2_dlygate4sd3_1
X_06090_ net2844 net3428 net956 _00266_ VPWR VGND sg13g2_mux2_1
XFILLER_7_261 VPWR VGND sg13g2_fill_2
Xhold217 i_exotiny._1160_\[1\] VPWR VGND net2044 sg13g2_dlygate4sd3_1
Xhold228 _03181_ VPWR VGND net2055 sg13g2_dlygate4sd3_1
X_08040__654 VPWR VGND net654 sg13g2_tiehi
X_05041_ net1238 net1240 _01768_ _01773_ VPWR VGND sg13g2_nor3_2
Xhold239 _01046_ VPWR VGND net2066 sg13g2_dlygate4sd3_1
X_08800_ net1608 VGND VPWR _00858_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[31\]
+ clknet_leaf_166_clk_regs sg13g2_dfrbpq_1
X_06992_ net2805 net875 _02922_ _02927_ VPWR VGND sg13g2_mux2_1
X_05943_ net2319 net2792 net968 _00152_ VPWR VGND sg13g2_mux2_1
XFILLER_67_942 VPWR VGND sg13g2_fill_2
X_08731_ net1677 VGND VPWR _00789_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[26\]
+ clknet_leaf_116_clk_regs sg13g2_dfrbpq_1
Xfanout1290 net1291 net1290 VPWR VGND sg13g2_buf_1
X_08662_ net775 VGND VPWR _00730_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[31\]
+ clknet_leaf_147_clk_regs sg13g2_dfrbpq_1
XFILLER_38_154 VPWR VGND sg13g2_fill_1
X_07613_ VGND VPWR i_exotiny.i_wdg_top.clk_div_inst.cnt\[15\] _03176_ _03179_ net1880
+ sg13g2_a21oi_1
XFILLER_93_282 VPWR VGND sg13g2_decap_8
XFILLER_54_636 VPWR VGND sg13g2_fill_1
X_05874_ net1184 _02460_ _02461_ VPWR VGND sg13g2_nor2_1
X_04825_ net1849 net1841 net1835 net1859 _01565_ VPWR VGND sg13g2_or4_1
X_08593_ net1803 VGND VPWR _00665_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data[0]
+ clknet_leaf_31_clk_regs sg13g2_dfrbpq_2
X_07544_ _03135_ net1883 net3586 VPWR VGND sg13g2_xnor2_1
X_04756_ VPWR VGND _01499_ net3694 _01478_ net1174 _01508_ _01454_ sg13g2_a221oi_1
X_04687_ i_exotiny._1489_\[0\] net1202 _01445_ net3523 net1266 VPWR VGND sg13g2_a22oi_1
X_07475_ net1211 net3825 _03018_ _01068_ VPWR VGND sg13g2_a21o_1
XFILLER_14_48 VPWR VGND sg13g2_fill_2
X_09214_ net765 VGND VPWR net2072 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[4\]
+ clknet_leaf_135_clk_regs sg13g2_dfrbpq_1
X_06426_ _01489_ _01513_ _02604_ VPWR VGND sg13g2_nor2_1
X_06357_ net3432 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[12\]
+ net1028 _00487_ VPWR VGND sg13g2_mux2_1
X_09145_ net837 VGND VPWR _01200_ i_exotiny._0027_\[1\] clknet_leaf_172_clk_regs sg13g2_dfrbpq_2
X_09076_ net1326 VGND VPWR net1882 i_exotiny.i_wdg_top.clk_div_inst.cnt\[16\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_06288_ net2778 net2698 net941 _00431_ VPWR VGND sg13g2_mux2_1
X_05308_ _02027_ _02028_ _02026_ _02034_ VPWR VGND _02033_ sg13g2_nand4_1
X_08027_ net667 VGND VPWR _00108_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[28\]
+ clknet_leaf_63_clk_regs sg13g2_dfrbpq_1
X_05239_ i_exotiny._0036_\[1\] _01644_ _01967_ VPWR VGND sg13g2_nor2_1
XFILLER_104_811 VPWR VGND sg13g2_decap_8
Xhold773 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[5\]
+ VPWR VGND net2600 sg13g2_dlygate4sd3_1
Xhold751 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[11\]
+ VPWR VGND net2578 sg13g2_dlygate4sd3_1
Xhold740 _00365_ VPWR VGND net2567 sg13g2_dlygate4sd3_1
Xhold762 _00245_ VPWR VGND net2589 sg13g2_dlygate4sd3_1
XFILLER_103_332 VPWR VGND sg13g2_decap_8
Xhold795 _00395_ VPWR VGND net2622 sg13g2_dlygate4sd3_1
Xhold784 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[11\]
+ VPWR VGND net2611 sg13g2_dlygate4sd3_1
XFILLER_104_888 VPWR VGND sg13g2_decap_8
X_09303__937 VPWR VGND net1357 sg13g2_tiehi
X_08929_ net1473 VGND VPWR _00987_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[27\]
+ clknet_leaf_65_clk_regs sg13g2_dfrbpq_1
Xhold1451 _00319_ VPWR VGND net3278 sg13g2_dlygate4sd3_1
Xhold1440 _00458_ VPWR VGND net3267 sg13g2_dlygate4sd3_1
Xhold1462 _00742_ VPWR VGND net3289 sg13g2_dlygate4sd3_1
Xhold1495 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[30\]
+ VPWR VGND net3322 sg13g2_dlygate4sd3_1
Xhold1484 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[17\]
+ VPWR VGND net3311 sg13g2_dlygate4sd3_1
Xhold1473 _00713_ VPWR VGND net3300 sg13g2_dlygate4sd3_1
XFILLER_44_113 VPWR VGND sg13g2_fill_2
X_08484__196 VPWR VGND net196 sg13g2_tiehi
XFILLER_44_157 VPWR VGND sg13g2_fill_1
XFILLER_71_65 VPWR VGND sg13g2_fill_1
XFILLER_9_515 VPWR VGND sg13g2_fill_2
XFILLER_40_352 VPWR VGND sg13g2_fill_1
XFILLER_41_875 VPWR VGND sg13g2_fill_2
XFILLER_40_385 VPWR VGND sg13g2_fill_2
XFILLER_41_897 VPWR VGND sg13g2_fill_2
X_08393__533 VPWR VGND net533 sg13g2_tiehi
Xclkbuf_leaf_120_clk_regs clknet_5_22__leaf_clk_regs clknet_leaf_120_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_5_776 VPWR VGND sg13g2_decap_8
XFILLER_106_181 VPWR VGND sg13g2_decap_8
X_08491__189 VPWR VGND net189 sg13g2_tiehi
X_08317__361 VPWR VGND net361 sg13g2_tiehi
XFILLER_1_971 VPWR VGND sg13g2_decap_8
X_08852__1134 VPWR VGND net1554 sg13g2_tiehi
XFILLER_64_945 VPWR VGND sg13g2_fill_2
XFILLER_64_967 VPWR VGND sg13g2_fill_1
X_04610_ VPWR _01372_ _00019_ VGND sg13g2_inv_1
XFILLER_51_628 VPWR VGND sg13g2_decap_8
X_05590_ i_exotiny._0352_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.carry_r
+ _02264_ VPWR VGND sg13g2_nor2_1
XFILLER_90_296 VPWR VGND sg13g2_fill_1
X_08324__354 VPWR VGND net354 sg13g2_tiehi
X_07260_ net2542 net2454 net1004 _00983_ VPWR VGND sg13g2_mux2_1
X_07191_ _02960_ net3606 net1111 VPWR VGND sg13g2_nand2_1
X_06211_ net2475 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[19\]
+ net949 _00366_ VPWR VGND sg13g2_mux2_1
X_08596__1380 VPWR VGND net1800 sg13g2_tiehi
X_06142_ _02528_ net3302 net1043 _00310_ VPWR VGND sg13g2_mux2_1
X_06073_ _02519_ net1139 net1166 _02520_ VPWR VGND sg13g2_a21o_2
X_05024_ _01756_ net1238 VPWR VGND net1240 sg13g2_nand2b_2
XFILLER_99_842 VPWR VGND sg13g2_decap_8
XFILLER_98_341 VPWR VGND sg13g2_decap_8
XFILLER_101_836 VPWR VGND sg13g2_decap_8
XFILLER_100_346 VPWR VGND sg13g2_decap_8
X_08331__347 VPWR VGND net347 sg13g2_tiehi
X_06975_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[17\]
+ net1994 net1018 _00748_ VPWR VGND sg13g2_mux2_1
X_08714_ net1694 VGND VPWR _00772_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[9\]
+ clknet_leaf_121_clk_regs sg13g2_dfrbpq_1
X_05926_ net2444 _02481_ net972 _00141_ VPWR VGND sg13g2_mux2_1
XFILLER_55_912 VPWR VGND sg13g2_fill_2
XFILLER_70_904 VPWR VGND sg13g2_fill_2
X_05857_ _02445_ net3306 net1053 _00108_ VPWR VGND sg13g2_mux2_1
X_08645_ net1752 VGND VPWR net3300 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[14\]
+ clknet_leaf_147_clk_regs sg13g2_dfrbpq_1
X_04808_ _01552_ VPWR _00009_ VGND _01485_ _01492_ sg13g2_o21ai_1
X_08576_ net52 VGND VPWR net2009 i_exotiny._0314_\[21\] clknet_leaf_181_clk_regs sg13g2_dfrbpq_1
X_05788_ net3792 VPWR _00075_ VGND _02390_ _02408_ sg13g2_o21ai_1
X_07527_ _01499_ _02471_ _03123_ VPWR VGND sg13g2_nor2_1
X_04739_ net3521 VPWR _00007_ VGND net1146 _01492_ sg13g2_o21ai_1
XFILLER_50_661 VPWR VGND sg13g2_decap_8
X_09190__791 VPWR VGND net791 sg13g2_tiehi
XFILLER_10_514 VPWR VGND sg13g2_fill_1
XFILLER_23_897 VPWR VGND sg13g2_fill_2
X_07458_ _03095_ net1148 _03032_ net1208 net1911 VPWR VGND sg13g2_a22oi_1
X_07389_ VGND VPWR net1078 _03042_ _01043_ _03040_ sg13g2_a21oi_1
XFILLER_41_57 VPWR VGND sg13g2_fill_2
X_06409_ VPWR VGND _02591_ _01553_ _02571_ _01520_ _02592_ _02226_ sg13g2_a221oi_1
X_09128_ net854 VGND VPWR _01183_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[16\]
+ clknet_leaf_152_clk_regs sg13g2_dfrbpq_1
X_08023__671 VPWR VGND net671 sg13g2_tiehi
X_09059_ net1343 VGND VPWR net3701 i_exotiny.i_wb_qspi_mem.cnt_r\[2\] clknet_leaf_27_clk_regs
+ sg13g2_dfrbpq_2
Xhold581 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[6\]
+ VPWR VGND net2408 sg13g2_dlygate4sd3_1
Xhold570 _01156_ VPWR VGND net2397 sg13g2_dlygate4sd3_1
Xhold592 _00149_ VPWR VGND net2419 sg13g2_dlygate4sd3_1
XFILLER_2_768 VPWR VGND sg13g2_decap_8
XFILLER_89_396 VPWR VGND sg13g2_fill_2
X_08633__1344 VPWR VGND net1764 sg13g2_tiehi
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_106_83 VPWR VGND sg13g2_decap_8
Xhold1270 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[29\]
+ VPWR VGND net3097 sg13g2_dlygate4sd3_1
Xhold1281 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[19\]
+ VPWR VGND net3108 sg13g2_dlygate4sd3_1
Xhold1292 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[8\]
+ VPWR VGND net3119 sg13g2_dlygate4sd3_1
XFILLER_82_31 VPWR VGND sg13g2_fill_2
XFILLER_46_989 VPWR VGND sg13g2_fill_2
X_08030__664 VPWR VGND net664 sg13g2_tiehi
XFILLER_61_959 VPWR VGND sg13g2_fill_1
XFILLER_14_831 VPWR VGND sg13g2_fill_2
XFILLER_60_458 VPWR VGND sg13g2_fill_1
XFILLER_9_301 VPWR VGND sg13g2_fill_1
XFILLER_13_330 VPWR VGND sg13g2_fill_1
XFILLER_95_300 VPWR VGND sg13g2_decap_8
XFILLER_68_525 VPWR VGND sg13g2_fill_2
XFILLER_83_528 VPWR VGND sg13g2_fill_2
X_06760_ _02786_ VPWR _02787_ VGND net3622 _02720_ sg13g2_o21ai_1
XFILLER_55_219 VPWR VGND sg13g2_fill_1
X_05711_ net1114 i_exotiny._1924_\[28\] _02354_ VPWR VGND sg13g2_nor2b_1
X_06691_ _02728_ net1187 net2014 VPWR VGND sg13g2_nand2b_1
X_08430_ net255 VGND VPWR net2577 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[29\]
+ clknet_leaf_91_clk_regs sg13g2_dfrbpq_1
X_05642_ VGND VPWR net1065 _02302_ _00036_ _02300_ sg13g2_a21oi_1
XFILLER_64_775 VPWR VGND sg13g2_fill_2
XFILLER_64_764 VPWR VGND sg13g2_fill_1
X_08788__1200 VPWR VGND net1620 sg13g2_tiehi
XFILLER_36_466 VPWR VGND sg13g2_fill_1
X_08361_ net317 VGND VPWR _00442_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[31\]
+ clknet_leaf_99_clk_regs sg13g2_dfrbpq_1
X_05573_ VGND VPWR net1202 _02250_ _02253_ _02252_ sg13g2_a21oi_1
X_08292_ net386 VGND VPWR _00373_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[26\]
+ clknet_leaf_106_clk_regs sg13g2_dfrbpq_1
X_07312_ net1253 net3798 net1150 _01024_ VPWR VGND sg13g2_mux2_1
X_07243_ net2361 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[6\]
+ net1003 _00966_ VPWR VGND sg13g2_mux2_1
XFILLER_31_182 VPWR VGND sg13g2_fill_2
X_08711__1277 VPWR VGND net1697 sg13g2_tiehi
X_07174_ _02950_ net2660 net1008 _00920_ VPWR VGND sg13g2_mux2_1
X_08007__688 VPWR VGND net688 sg13g2_tiehi
X_06125_ net3014 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[12\]
+ net1043 _00294_ VPWR VGND sg13g2_mux2_1
XFILLER_105_438 VPWR VGND sg13g2_decap_8
X_06056_ net2588 net2257 net964 _00241_ VPWR VGND sg13g2_mux2_1
XFILLER_87_801 VPWR VGND sg13g2_fill_1
X_05007_ _01738_ _01722_ _01701_ _01739_ VPWR VGND sg13g2_a21o_2
X_08933__1049 VPWR VGND net1469 sg13g2_tiehi
X_06958_ net2450 net3436 net1021 _00731_ VPWR VGND sg13g2_mux2_1
X_05909_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[14\]
+ net2351 net974 _00126_ VPWR VGND sg13g2_mux2_1
X_09077__905 VPWR VGND net1325 sg13g2_tiehi
X_06889_ net1128 _02893_ _02894_ _02895_ VPWR VGND sg13g2_nor3_1
XFILLER_15_617 VPWR VGND sg13g2_fill_2
X_08628_ net743 VGND VPWR net3679 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[1\]
+ clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
XFILLER_28_989 VPWR VGND sg13g2_fill_2
X_09255__552 VPWR VGND net552 sg13g2_tiehi
X_08559_ net92 VGND VPWR net3477 i_exotiny._0314_\[4\] clknet_leaf_181_clk_regs sg13g2_dfrbpq_1
X_08481__199 VPWR VGND net199 sg13g2_tiehi
X_08307__371 VPWR VGND net371 sg13g2_tiehi
XFILLER_7_805 VPWR VGND sg13g2_fill_2
XFILLER_105_972 VPWR VGND sg13g2_decap_8
XFILLER_104_460 VPWR VGND sg13g2_decap_8
X_08314__364 VPWR VGND net364 sg13g2_tiehi
XFILLER_92_314 VPWR VGND sg13g2_fill_1
Xfanout880 _02463_ net880 VPWR VGND sg13g2_buf_8
Xfanout891 net892 net891 VPWR VGND sg13g2_buf_8
X_08909__1073 VPWR VGND net1493 sg13g2_tiehi
XFILLER_61_767 VPWR VGND sg13g2_fill_1
XFILLER_9_131 VPWR VGND sg13g2_fill_1
X_08321__357 VPWR VGND net357 sg13g2_tiehi
XFILLER_6_871 VPWR VGND sg13g2_decap_8
XFILLER_103_909 VPWR VGND sg13g2_decap_8
X_07930_ net718 VGND VPWR net2047 i_exotiny._1924_\[23\] clknet_leaf_25_clk_regs sg13g2_dfrbpq_1
X_07861_ _03228_ net1142 net1163 _03229_ VPWR VGND sg13g2_a21o_2
X_06812_ VGND VPWR net3563 net1132 _02831_ _02830_ sg13g2_a21oi_1
XFILLER_3_1012 VPWR VGND sg13g2_decap_8
X_07792_ net3481 net3323 net894 _01271_ VPWR VGND sg13g2_mux2_1
X_06743_ VGND VPWR net1101 _02771_ _00667_ _02772_ sg13g2_a21oi_1
X_08729__1259 VPWR VGND net1679 sg13g2_tiehi
X_06674_ VPWR VGND _02711_ net1195 _02710_ _01369_ _00659_ net1153 sg13g2_a221oi_1
X_08413_ net272 VGND VPWR net3433 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[12\]
+ clknet_leaf_91_clk_regs sg13g2_dfrbpq_1
X_08013__681 VPWR VGND net681 sg13g2_tiehi
X_05625_ VGND VPWR i_exotiny._1612_\[2\] net1124 _02290_ _02289_ sg13g2_a21oi_1
X_08344_ net334 VGND VPWR _00425_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[14\]
+ clknet_leaf_95_clk_regs sg13g2_dfrbpq_1
X_05556_ net1277 i_exotiny._0315_\[22\] _02239_ VPWR VGND sg13g2_nor2b_1
X_08275_ net403 VGND VPWR _00356_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[9\]
+ clknet_leaf_99_clk_regs sg13g2_dfrbpq_1
X_05487_ _02185_ net3457 net1069 VPWR VGND sg13g2_nand2_1
X_07226_ net3587 i_exotiny.i_wb_spi.dat_rx_r\[23\] net1087 _00951_ VPWR VGND sg13g2_mux2_1
X_07157_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[18\]
+ net3214 net1010 _00905_ VPWR VGND sg13g2_mux2_1
XFILLER_105_235 VPWR VGND sg13g2_decap_8
X_06108_ net3412 net874 _02519_ _02524_ VPWR VGND sg13g2_mux2_1
XFILLER_106_769 VPWR VGND sg13g2_decap_8
X_07088_ net2967 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[20\]
+ net913 _00843_ VPWR VGND sg13g2_mux2_1
X_08020__674 VPWR VGND net674 sg13g2_tiehi
Xfanout1119 net1120 net1119 VPWR VGND sg13g2_buf_8
X_06039_ net2611 net2513 net963 _00224_ VPWR VGND sg13g2_mux2_1
Xfanout1108 _01686_ net1108 VPWR VGND sg13g2_buf_2
XFILLER_59_333 VPWR VGND sg13g2_fill_1
XFILLER_102_986 VPWR VGND sg13g2_decap_8
XFILLER_101_485 VPWR VGND sg13g2_decap_8
XFILLER_90_829 VPWR VGND sg13g2_fill_1
XFILLER_103_62 VPWR VGND sg13g2_fill_1
XFILLER_43_734 VPWR VGND sg13g2_fill_2
XFILLER_11_642 VPWR VGND sg13g2_fill_1
XFILLER_42_299 VPWR VGND sg13g2_fill_2
XFILLER_10_163 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_98_clk_regs clknet_5_29__leaf_clk_regs clknet_leaf_98_clk_regs VPWR VGND
+ sg13g2_buf_8
Xclkbuf_leaf_27_clk_regs clknet_5_9__leaf_clk_regs clknet_leaf_27_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_3_830 VPWR VGND sg13g2_decap_8
XFILLER_40_9 VPWR VGND sg13g2_fill_2
XFILLER_92_100 VPWR VGND sg13g2_fill_1
XFILLER_81_818 VPWR VGND sg13g2_fill_2
X_05410_ net1113 _02120_ _02121_ i_exotiny._2043_\[7\] VPWR VGND sg13g2_nor3_1
XFILLER_33_255 VPWR VGND sg13g2_fill_2
XFILLER_15_992 VPWR VGND sg13g2_fill_1
X_06390_ _02577_ net3493 net1271 VPWR VGND sg13g2_nand2_1
X_05341_ VGND VPWR _02065_ _02064_ _02063_ sg13g2_or2_1
XFILLER_88_1007 VPWR VGND sg13g2_decap_8
X_08060_ net634 VGND VPWR net2445 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[29\]
+ clknet_leaf_55_clk_regs sg13g2_dfrbpq_1
X_05272_ _01998_ _01791_ i_exotiny._0026_\[0\] _01758_ i_exotiny._0040_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_07011_ net3130 net2912 net918 _00778_ VPWR VGND sg13g2_mux2_1
X_09067__915 VPWR VGND net1335 sg13g2_tiehi
XFILLER_52_0 VPWR VGND sg13g2_decap_8
X_08962_ net1440 VGND VPWR net3233 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[28\]
+ clknet_leaf_75_clk_regs sg13g2_dfrbpq_1
X_09245__562 VPWR VGND net562 sg13g2_tiehi
XFILLER_102_238 VPWR VGND sg13g2_decap_8
XFILLER_97_940 VPWR VGND sg13g2_decap_8
X_07913_ net735 VGND VPWR net1988 i_exotiny._1924_\[6\] clknet_leaf_33_clk_regs sg13g2_dfrbpq_1
X_08893_ net1509 VGND VPWR net3588 i_exotiny.i_wb_spi.dat_rx_r\[23\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_96_472 VPWR VGND sg13g2_decap_4
Xhold1803 i_exotiny._1614_\[2\] VPWR VGND net3630 sg13g2_dlygate4sd3_1
Xhold1836 i_exotiny.i_wb_spi.dat_rx_r\[24\] VPWR VGND net3663 sg13g2_dlygate4sd3_1
Xhold1825 _01547_ VPWR VGND net3652 sg13g2_dlygate4sd3_1
Xhold1814 i_exotiny._0369_\[11\] VPWR VGND net3641 sg13g2_dlygate4sd3_1
X_07844_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[24\]
+ net2469 net986 _01317_ VPWR VGND sg13g2_mux2_1
Xhold1847 i_exotiny._0014_\[2\] VPWR VGND net3674 sg13g2_dlygate4sd3_1
Xhold1869 _00005_ VPWR VGND net3696 sg13g2_dlygate4sd3_1
Xhold1858 _01028_ VPWR VGND net3685 sg13g2_dlygate4sd3_1
X_07775_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[31\]
+ net2559 net990 _01260_ VPWR VGND sg13g2_mux2_1
X_08571__62 VPWR VGND net62 sg13g2_tiehi
X_04987_ _01712_ _01718_ _01719_ VPWR VGND sg13g2_nor2_1
X_06726_ net1173 VPWR _02758_ VGND i_exotiny._0369_\[5\] net1193 sg13g2_o21ai_1
X_09074__908 VPWR VGND net1328 sg13g2_tiehi
XFILLER_80_862 VPWR VGND sg13g2_fill_2
X_06657_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.carry_r[0] i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[0\].i_hadd.a_i
+ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[1\].i_hadd.a_i _02697_
+ VPWR VGND sg13g2_a21o_1
X_05608_ VGND VPWR i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_sw_write_data[0]
+ net1118 _02277_ _02276_ sg13g2_a21oi_1
X_08865__1121 VPWR VGND net1541 sg13g2_tiehi
XFILLER_52_575 VPWR VGND sg13g2_fill_1
XFILLER_25_778 VPWR VGND sg13g2_fill_1
X_09252__555 VPWR VGND net555 sg13g2_tiehi
X_06588_ net1194 _02647_ _02648_ _00636_ VPWR VGND sg13g2_nor3_1
X_08327_ net351 VGND VPWR net3165 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[29\]
+ clknet_leaf_72_clk_regs sg13g2_dfrbpq_1
X_08883__1099 VPWR VGND net1519 sg13g2_tiehi
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
X_05539_ i_exotiny.i_wb_qspi_mem.crm_r net1218 _02226_ VPWR VGND sg13g2_nor2_1
X_08304__374 VPWR VGND net374 sg13g2_tiehi
X_08258_ net419 VGND VPWR _00339_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[25\]
+ clknet_leaf_57_clk_regs sg13g2_dfrbpq_1
XFILLER_20_483 VPWR VGND sg13g2_fill_1
X_07209_ net1897 net1089 _02966_ VPWR VGND sg13g2_nor2_1
X_08189_ net488 VGND VPWR net2799 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[20\]
+ clknet_leaf_110_clk_regs sg13g2_dfrbpq_1
XFILLER_106_566 VPWR VGND sg13g2_decap_8
XFILLER_88_951 VPWR VGND sg13g2_decap_8
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_102_783 VPWR VGND sg13g2_decap_8
XFILLER_101_282 VPWR VGND sg13g2_decap_8
X_08311__367 VPWR VGND net367 sg13g2_tiehi
XFILLER_74_155 VPWR VGND sg13g2_fill_2
XFILLER_74_144 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_145_clk_regs clknet_5_16__leaf_clk_regs clknet_leaf_145_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_74_177 VPWR VGND sg13g2_fill_1
XFILLER_56_892 VPWR VGND sg13g2_fill_2
X_07904__43 VPWR VGND net43 sg13g2_tiehi
XFILLER_15_266 VPWR VGND sg13g2_fill_2
XFILLER_43_564 VPWR VGND sg13g2_fill_1
XFILLER_8_944 VPWR VGND sg13g2_decap_8
X_09275__71 VPWR VGND net71 sg13g2_tiehi
XFILLER_12_995 VPWR VGND sg13g2_decap_8
XFILLER_3_660 VPWR VGND sg13g2_fill_2
X_04910_ net1258 net1261 net1256 _01642_ VGND VPWR _01640_ sg13g2_nor4_2
X_05890_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[1\] _02474_ _02475_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_94_976 VPWR VGND sg13g2_decap_8
X_04841_ net1111 _01580_ _01581_ VPWR VGND sg13g2_nor2_1
XFILLER_19_550 VPWR VGND sg13g2_fill_1
XFILLER_94_1011 VPWR VGND sg13g2_decap_8
X_07560_ net3833 net3520 net3724 _01521_ _03145_ VPWR VGND sg13g2_nor4_1
XFILLER_0_1015 VPWR VGND sg13g2_decap_8
X_04772_ _01513_ VPWR _01523_ VGND _01521_ _01522_ sg13g2_o21ai_1
X_06511_ net3031 net2835 net932 _00586_ VPWR VGND sg13g2_mux2_1
X_08646__1331 VPWR VGND net1751 sg13g2_tiehi
X_09230_ net749 VGND VPWR net3226 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[20\]
+ clknet_leaf_136_clk_regs sg13g2_dfrbpq_1
X_07491_ VGND VPWR _01393_ net906 _01075_ _03112_ sg13g2_a21oi_1
X_06442_ net2057 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[7\]
+ net934 _00529_ VPWR VGND sg13g2_mux2_1
X_06373_ i_exotiny._0035_\[0\] net889 _02565_ _02567_ VPWR VGND sg13g2_mux2_1
X_09161_ net821 VGND VPWR _01216_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[17\]
+ clknet_leaf_173_clk_regs sg13g2_dfrbpq_1
XFILLER_21_258 VPWR VGND sg13g2_fill_2
X_08112_ net582 VGND VPWR net3488 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[17\]
+ clknet_leaf_124_clk_regs sg13g2_dfrbpq_1
X_09092_ net1310 VGND VPWR _01147_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[12\]
+ clknet_leaf_141_clk_regs sg13g2_dfrbpq_1
X_05324_ _02041_ _02045_ _02046_ _02048_ VPWR VGND sg13g2_nor3_1
X_08043_ net651 VGND VPWR _00124_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[12\]
+ clknet_leaf_53_clk_regs sg13g2_dfrbpq_1
Xhold911 _00538_ VPWR VGND net2738 sg13g2_dlygate4sd3_1
Xhold922 _01220_ VPWR VGND net2749 sg13g2_dlygate4sd3_1
Xhold900 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[29\]
+ VPWR VGND net2727 sg13g2_dlygate4sd3_1
X_05255_ VGND VPWR _01981_ _01742_ _01715_ sg13g2_or2_1
Xhold944 _00753_ VPWR VGND net2771 sg13g2_dlygate4sd3_1
Xhold933 _00984_ VPWR VGND net2760 sg13g2_dlygate4sd3_1
Xhold955 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[27\]
+ VPWR VGND net2782 sg13g2_dlygate4sd3_1
X_05186_ VGND VPWR _01743_ _01913_ _01914_ _01702_ sg13g2_a21oi_1
XFILLER_103_514 VPWR VGND sg13g2_decap_8
Xhold966 _00156_ VPWR VGND net2793 sg13g2_dlygate4sd3_1
Xhold988 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[5\]
+ VPWR VGND net2815 sg13g2_dlygate4sd3_1
Xhold977 i_exotiny._0021_\[3\] VPWR VGND net2804 sg13g2_dlygate4sd3_1
Xhold999 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[11\]
+ VPWR VGND net2826 sg13g2_dlygate4sd3_1
X_08945_ net1457 VGND VPWR net2790 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[11\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
XFILLER_69_461 VPWR VGND sg13g2_decap_4
Xhold1600 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[22\]
+ VPWR VGND net3427 sg13g2_dlygate4sd3_1
Xhold1622 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[11\]
+ VPWR VGND net3449 sg13g2_dlygate4sd3_1
Xhold1644 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[27\]
+ VPWR VGND net3471 sg13g2_dlygate4sd3_1
XFILLER_96_280 VPWR VGND sg13g2_decap_8
Xhold1633 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[13\]
+ VPWR VGND net3460 sg13g2_dlygate4sd3_1
X_08876_ net1526 VGND VPWR _00934_ i_exotiny.i_wb_spi.dat_rx_r\[6\] clknet_leaf_24_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_57_645 VPWR VGND sg13g2_fill_1
X_08119__575 VPWR VGND net575 sg13g2_tiehi
Xhold1611 _00922_ VPWR VGND net3438 sg13g2_dlygate4sd3_1
Xhold1655 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[6\]
+ VPWR VGND net3482 sg13g2_dlygate4sd3_1
Xhold1666 i_exotiny._0314_\[4\] VPWR VGND net3493 sg13g2_dlygate4sd3_1
Xhold1677 i_exotiny._0314_\[13\] VPWR VGND net3504 sg13g2_dlygate4sd3_1
X_07827_ net2307 i_exotiny._0022_\[3\] net984 _01300_ VPWR VGND sg13g2_mux2_1
X_07758_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[14\]
+ net3057 net988 _01243_ VPWR VGND sg13g2_mux2_1
Xhold1688 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[5\]
+ VPWR VGND net3515 sg13g2_dlygate4sd3_1
XFILLER_57_689 VPWR VGND sg13g2_fill_1
Xhold1699 i_exotiny._1160_\[11\] VPWR VGND net3526 sg13g2_dlygate4sd3_1
X_06709_ VPWR VGND _02742_ _02741_ net1173 net3666 _02744_ net1181 sg13g2_a221oi_1
XFILLER_71_169 VPWR VGND sg13g2_fill_1
XFILLER_13_704 VPWR VGND sg13g2_fill_1
X_07689_ net2526 net2976 net1000 _01191_ VPWR VGND sg13g2_mux2_1
XFILLER_44_46 VPWR VGND sg13g2_fill_1
XFILLER_52_372 VPWR VGND sg13g2_fill_2
X_08126__568 VPWR VGND net568 sg13g2_tiehi
XFILLER_5_903 VPWR VGND sg13g2_decap_8
XFILLER_20_280 VPWR VGND sg13g2_fill_2
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_4_413 VPWR VGND sg13g2_fill_1
XFILLER_106_363 VPWR VGND sg13g2_decap_8
XFILLER_79_214 VPWR VGND sg13g2_fill_1
XFILLER_4_479 VPWR VGND sg13g2_fill_1
X_08724__1264 VPWR VGND net1684 sg13g2_tiehi
XFILLER_0_663 VPWR VGND sg13g2_fill_2
XFILLER_47_111 VPWR VGND sg13g2_fill_1
XFILLER_78_1028 VPWR VGND sg13g2_fill_1
X_09057__925 VPWR VGND net1345 sg13g2_tiehi
X_08946__1036 VPWR VGND net1456 sg13g2_tiehi
XFILLER_16_597 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_42_clk_regs clknet_5_10__leaf_clk_regs clknet_leaf_42_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_15_1023 VPWR VGND sg13g2_decap_4
Xhold207 _00058_ VPWR VGND net2034 sg13g2_dlygate4sd3_1
Xhold229 _01132_ VPWR VGND net2056 sg13g2_dlygate4sd3_1
X_05040_ net1220 _01754_ _01762_ _01772_ VPWR VGND sg13g2_nor3_2
Xhold218 _01038_ VPWR VGND net2045 sg13g2_dlygate4sd3_1
X_09064__918 VPWR VGND net1338 sg13g2_tiehi
XFILLER_98_523 VPWR VGND sg13g2_fill_2
X_06991_ net2160 _02926_ net1020 _00761_ VPWR VGND sg13g2_mux2_1
X_09242__565 VPWR VGND net565 sg13g2_tiehi
XFILLER_100_528 VPWR VGND sg13g2_decap_8
X_05942_ net3081 net3378 net966 _00151_ VPWR VGND sg13g2_mux2_1
X_08730_ net1678 VGND VPWR _00788_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[25\]
+ clknet_leaf_121_clk_regs sg13g2_dfrbpq_1
Xfanout1291 net3571 net1291 VPWR VGND sg13g2_buf_8
X_08661_ net1736 VGND VPWR _00729_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[30\]
+ clknet_leaf_149_clk_regs sg13g2_dfrbpq_1
XFILLER_22_1027 VPWR VGND sg13g2_fill_2
X_05873_ _02429_ _02459_ _02460_ VPWR VGND sg13g2_nor2_1
Xfanout1280 i_exotiny._1312_ net1280 VPWR VGND sg13g2_buf_2
X_07612_ net1205 net3650 _01130_ VPWR VGND sg13g2_nor2_1
X_04824_ _01561_ _01563_ _01560_ _01564_ VPWR VGND sg13g2_nand3_1
XFILLER_26_306 VPWR VGND sg13g2_fill_1
XFILLER_39_689 VPWR VGND sg13g2_fill_1
X_08592_ net1804 VGND VPWR _00664_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data[0]
+ clknet_leaf_28_clk_regs sg13g2_dfrbpq_2
X_07543_ net1883 _03133_ _01105_ VPWR VGND sg13g2_nor2_1
XFILLER_41_309 VPWR VGND sg13g2_fill_1
X_04755_ _01507_ net1174 _01454_ VPWR VGND sg13g2_nand2_2
X_04686_ net1266 i_exotiny._0315_\[6\] _01445_ VPWR VGND sg13g2_nor2_1
X_07474_ net1211 net3826 _03083_ _01067_ VPWR VGND sg13g2_a21o_1
X_06425_ _00518_ _02602_ _02603_ VPWR VGND sg13g2_nand2_1
X_09213_ net766 VGND VPWR _01268_ i_exotiny._0023_\[3\] clknet_leaf_130_clk_regs sg13g2_dfrbpq_2
X_08802__1186 VPWR VGND net1606 sg13g2_tiehi
X_09144_ net838 VGND VPWR net2993 i_exotiny._0027_\[0\] clknet_leaf_174_clk_regs sg13g2_dfrbpq_2
X_06356_ net2851 net2269 net1030 _00486_ VPWR VGND sg13g2_mux2_1
X_09075_ net1327 VGND VPWR _01130_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[15\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_06287_ net2820 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[19\]
+ net943 _00430_ VPWR VGND sg13g2_mux2_1
X_05307_ _02029_ _02030_ _02031_ _02032_ _02033_ VPWR VGND sg13g2_and4_1
Xhold730 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[10\]
+ VPWR VGND net2557 sg13g2_dlygate4sd3_1
X_08301__377 VPWR VGND net377 sg13g2_tiehi
X_08026_ net668 VGND VPWR net2092 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[27\]
+ clknet_leaf_59_clk_regs sg13g2_dfrbpq_1
X_05238_ _01950_ _01955_ _01965_ _01966_ VPWR VGND sg13g2_nor3_2
XFILLER_89_501 VPWR VGND sg13g2_fill_1
Xhold763 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[11\]
+ VPWR VGND net2590 sg13g2_dlygate4sd3_1
Xhold752 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[13\]
+ VPWR VGND net2579 sg13g2_dlygate4sd3_1
Xhold741 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[19\]
+ VPWR VGND net2568 sg13g2_dlygate4sd3_1
XFILLER_104_867 VPWR VGND sg13g2_decap_8
XFILLER_103_311 VPWR VGND sg13g2_decap_8
Xhold774 _01234_ VPWR VGND net2601 sg13g2_dlygate4sd3_1
Xhold796 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[25\]
+ VPWR VGND net2623 sg13g2_dlygate4sd3_1
Xhold785 _00228_ VPWR VGND net2612 sg13g2_dlygate4sd3_1
X_05169_ net1110 _01897_ _01899_ VPWR VGND sg13g2_and2_1
XFILLER_103_388 VPWR VGND sg13g2_decap_8
X_08928_ net1474 VGND VPWR _00986_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[26\]
+ clknet_leaf_19_clk_regs sg13g2_dfrbpq_1
Xhold1452 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[21\]
+ VPWR VGND net3279 sg13g2_dlygate4sd3_1
Xhold1430 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[14\]
+ VPWR VGND net3257 sg13g2_dlygate4sd3_1
Xhold1441 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[10\]
+ VPWR VGND net3268 sg13g2_dlygate4sd3_1
XFILLER_29_133 VPWR VGND sg13g2_fill_1
Xhold1463 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[24\]
+ VPWR VGND net3290 sg13g2_dlygate4sd3_1
XFILLER_85_773 VPWR VGND sg13g2_fill_2
Xhold1485 _01152_ VPWR VGND net3312 sg13g2_dlygate4sd3_1
X_08859_ net1547 VGND VPWR _00917_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[26\]
+ clknet_leaf_186_clk_regs sg13g2_dfrbpq_1
Xhold1474 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[31\]
+ VPWR VGND net3301 sg13g2_dlygate4sd3_1
Xhold1496 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[10\]
+ VPWR VGND net3323 sg13g2_dlygate4sd3_1
XFILLER_106_160 VPWR VGND sg13g2_decap_8
XFILLER_84_1010 VPWR VGND sg13g2_decap_8
XFILLER_1_950 VPWR VGND sg13g2_decap_8
XFILLER_45_1027 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_160_clk_regs clknet_5_7__leaf_clk_regs clknet_leaf_160_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_75_272 VPWR VGND sg13g2_fill_2
XFILLER_75_261 VPWR VGND sg13g2_fill_2
Xhold90 _00046_ VPWR VGND net1917 sg13g2_dlygate4sd3_1
XFILLER_36_604 VPWR VGND sg13g2_fill_2
XFILLER_91_776 VPWR VGND sg13g2_fill_1
XFILLER_90_275 VPWR VGND sg13g2_fill_2
X_06210_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[22\]
+ net2566 net948 _00365_ VPWR VGND sg13g2_mux2_1
XFILLER_32_898 VPWR VGND sg13g2_fill_1
X_07190_ VGND VPWR _01365_ _02956_ _00927_ net3745 sg13g2_a21oi_1
X_08109__585 VPWR VGND net585 sg13g2_tiehi
X_06141_ i_exotiny._0037_\[0\] net887 _02526_ _02528_ VPWR VGND sg13g2_mux2_1
X_06072_ _02517_ _02518_ _02519_ VPWR VGND sg13g2_nor2_2
XFILLER_99_821 VPWR VGND sg13g2_decap_8
X_05023_ net1221 _01753_ _01754_ _01755_ VPWR VGND sg13g2_or3_1
XFILLER_98_320 VPWR VGND sg13g2_decap_8
XFILLER_101_815 VPWR VGND sg13g2_decap_8
XFILLER_99_898 VPWR VGND sg13g2_decap_8
XFILLER_100_325 VPWR VGND sg13g2_decap_8
XFILLER_98_397 VPWR VGND sg13g2_decap_8
X_06974_ net2722 net2908 net1021 _00747_ VPWR VGND sg13g2_mux2_1
X_09179__802 VPWR VGND net802 sg13g2_tiehi
X_05925_ net881 i_exotiny._0019_\[1\] _02478_ _02481_ VPWR VGND sg13g2_mux2_1
X_08713_ net1695 VGND VPWR _00771_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[8\]
+ clknet_leaf_120_clk_regs sg13g2_dfrbpq_1
XFILLER_82_710 VPWR VGND sg13g2_fill_2
X_08116__578 VPWR VGND net578 sg13g2_tiehi
X_05856_ net3411 net886 _02421_ _02445_ VPWR VGND sg13g2_mux2_1
XFILLER_55_957 VPWR VGND sg13g2_fill_1
X_08644_ net1753 VGND VPWR net2266 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[13\]
+ clknet_leaf_147_clk_regs sg13g2_dfrbpq_1
X_05787_ _02409_ _01550_ _01372_ _01549_ net3791 VPWR VGND sg13g2_a22oi_1
X_04807_ _01552_ _01540_ _01541_ VPWR VGND sg13g2_nand2b_1
X_08575_ net54 VGND VPWR net2039 i_exotiny._0314_\[20\] clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
XFILLER_81_286 VPWR VGND sg13g2_fill_1
X_04738_ net3520 _01493_ net1283 _01494_ VPWR VGND sg13g2_nand3_1
X_07526_ _03122_ net2024 net901 VPWR VGND sg13g2_nand2_1
XFILLER_41_106 VPWR VGND sg13g2_decap_4
XFILLER_34_191 VPWR VGND sg13g2_fill_1
X_07457_ _03094_ net1911 net1212 VPWR VGND sg13g2_nand2_1
X_04669_ _01428_ _01429_ _01430_ VPWR VGND sg13g2_and2_1
X_06408_ i_exotiny._0315_\[20\] i_exotiny._0314_\[20\] net1271 _02591_ VPWR VGND sg13g2_mux2_1
X_07388_ _03042_ _03025_ _03041_ net1207 i_exotiny._1160_\[10\] VPWR VGND sg13g2_a22oi_1
X_06339_ _02562_ net2353 net1036 _00473_ VPWR VGND sg13g2_mux2_1
X_09127_ net855 VGND VPWR _01182_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[15\]
+ clknet_leaf_155_clk_regs sg13g2_dfrbpq_1
X_09058_ net1344 VGND VPWR net3725 i_exotiny.i_wb_qspi_mem.cnt_r\[1\] clknet_leaf_27_clk_regs
+ sg13g2_dfrbpq_2
X_08009_ net686 VGND VPWR net2599 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[10\]
+ clknet_leaf_68_clk_regs sg13g2_dfrbpq_1
Xhold571 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[29\]
+ VPWR VGND net2398 sg13g2_dlygate4sd3_1
Xhold560 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[27\]
+ VPWR VGND net2387 sg13g2_dlygate4sd3_1
XFILLER_2_747 VPWR VGND sg13g2_decap_8
XFILLER_104_664 VPWR VGND sg13g2_decap_8
X_08490__190 VPWR VGND net190 sg13g2_tiehi
Xhold582 _00701_ VPWR VGND net2409 sg13g2_dlygate4sd3_1
Xhold593 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[16\]
+ VPWR VGND net2420 sg13g2_dlygate4sd3_1
XFILLER_106_62 VPWR VGND sg13g2_decap_8
XFILLER_103_185 VPWR VGND sg13g2_decap_8
XFILLER_92_507 VPWR VGND sg13g2_fill_1
Xhold1260 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[10\]
+ VPWR VGND net3087 sg13g2_dlygate4sd3_1
XFILLER_66_55 VPWR VGND sg13g2_fill_1
Xhold1282 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[7\]
+ VPWR VGND net3109 sg13g2_dlygate4sd3_1
Xhold1293 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[28\]
+ VPWR VGND net3120 sg13g2_dlygate4sd3_1
Xhold1271 _01358_ VPWR VGND net3098 sg13g2_dlygate4sd3_1
XFILLER_60_404 VPWR VGND sg13g2_fill_1
XFILLER_54_990 VPWR VGND sg13g2_fill_1
X_09054__928 VPWR VGND net1348 sg13g2_tiehi
XFILLER_25_191 VPWR VGND sg13g2_fill_2
X_07985__126 VPWR VGND net126 sg13g2_tiehi
XFILLER_41_640 VPWR VGND sg13g2_fill_1
X_08896__1086 VPWR VGND net1506 sg13g2_tiehi
XFILLER_96_879 VPWR VGND sg13g2_decap_8
XFILLER_95_356 VPWR VGND sg13g2_decap_8
XFILLER_68_559 VPWR VGND sg13g2_fill_1
X_05710_ VGND VPWR net1058 _02353_ _00053_ _02351_ sg13g2_a21oi_1
X_06690_ VGND VPWR _02724_ _02726_ _02727_ _02721_ sg13g2_a21oi_1
X_05641_ VGND VPWR i_exotiny._1615_\[2\] net1124 _02302_ _02301_ sg13g2_a21oi_1
X_08360_ net318 VGND VPWR _00441_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[30\]
+ clknet_leaf_108_clk_regs sg13g2_dfrbpq_1
X_07311_ _02984_ net1212 net1196 VPWR VGND sg13g2_nand2b_1
X_05572_ net1201 _02251_ _02252_ VPWR VGND sg13g2_nor2_1
X_08291_ net387 VGND VPWR net2306 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[25\]
+ clknet_leaf_106_clk_regs sg13g2_dfrbpq_1
X_08683__1305 VPWR VGND net1725 sg13g2_tiehi
X_07242_ net2934 net2889 net1005 _00965_ VPWR VGND sg13g2_mux2_1
X_07173_ i_exotiny._0036_\[1\] net881 _02947_ _02950_ VPWR VGND sg13g2_mux2_1
X_06124_ net2602 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[11\]
+ net1044 _00293_ VPWR VGND sg13g2_mux2_1
XFILLER_105_417 VPWR VGND sg13g2_decap_8
X_06055_ net2657 net2018 net963 _00240_ VPWR VGND sg13g2_mux2_1
X_05006_ _01737_ _01730_ _01717_ _01738_ VPWR VGND sg13g2_a21o_1
X_08941__1041 VPWR VGND net1461 sg13g2_tiehi
XFILLER_74_507 VPWR VGND sg13g2_fill_2
X_06957_ _02922_ net1140 net1167 _02923_ VPWR VGND sg13g2_a21o_2
X_05908_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[13\]
+ net2883 net972 _00125_ VPWR VGND sg13g2_mux2_1
X_06888_ net1172 VPWR _02894_ VGND net3530 net1186 sg13g2_o21ai_1
XFILLER_55_754 VPWR VGND sg13g2_fill_1
X_08627_ net742 VGND VPWR net3524 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.macro_steps_r\[0\]
+ clknet_leaf_6_clk_regs sg13g2_dfrbpq_2
X_05839_ _01610_ _02425_ _02426_ _02427_ _02428_ VPWR VGND sg13g2_and4_1
XFILLER_54_297 VPWR VGND sg13g2_fill_1
XFILLER_52_13 VPWR VGND sg13g2_fill_2
XFILLER_23_651 VPWR VGND sg13g2_fill_1
X_08558_ net96 VGND VPWR _00631_ i_exotiny._0314_\[3\] clknet_leaf_5_clk_regs sg13g2_dfrbpq_2
X_08489_ net191 VGND VPWR net3020 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[9\]
+ clknet_leaf_70_clk_regs sg13g2_dfrbpq_1
X_07509_ net3113 i_exotiny._0315_\[22\] net905 _01092_ VPWR VGND sg13g2_mux2_1
XFILLER_50_492 VPWR VGND sg13g2_fill_2
XFILLER_10_345 VPWR VGND sg13g2_fill_2
XFILLER_105_951 VPWR VGND sg13g2_decap_8
Xhold390 _00854_ VPWR VGND net2217 sg13g2_dlygate4sd3_1
Xfanout881 net885 net881 VPWR VGND sg13g2_buf_8
Xfanout892 _03217_ net892 VPWR VGND sg13g2_buf_8
X_08761__1227 VPWR VGND net1647 sg13g2_tiehi
Xhold1090 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[7\]
+ VPWR VGND net2917 sg13g2_dlygate4sd3_1
XFILLER_18_467 VPWR VGND sg13g2_fill_1
XFILLER_45_231 VPWR VGND sg13g2_fill_1
XFILLER_60_234 VPWR VGND sg13g2_fill_2
XFILLER_14_651 VPWR VGND sg13g2_fill_1
XFILLER_9_187 VPWR VGND sg13g2_fill_2
XFILLER_6_850 VPWR VGND sg13g2_decap_8
X_08106__588 VPWR VGND net588 sg13g2_tiehi
XFILLER_54_4 VPWR VGND sg13g2_fill_1
XFILLER_69_802 VPWR VGND sg13g2_fill_1
X_07860_ _02477_ _02492_ _03228_ VPWR VGND sg13g2_nor2_2
X_06811_ net1132 _02828_ _02829_ _02830_ VPWR VGND sg13g2_nor3_1
X_07791_ net3203 net2833 net894 _01270_ VPWR VGND sg13g2_mux2_1
XFILLER_95_186 VPWR VGND sg13g2_fill_1
X_06742_ net3611 net1096 _02772_ VPWR VGND sg13g2_nor2_1
X_08737__1251 VPWR VGND net1671 sg13g2_tiehi
X_06673_ VGND VPWR net3611 _02690_ _02711_ net1153 sg13g2_a21oi_1
X_08412_ net273 VGND VPWR _00486_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[11\]
+ clknet_leaf_97_clk_regs sg13g2_dfrbpq_1
X_05624_ net1125 i_exotiny._1924_\[6\] _02289_ VPWR VGND sg13g2_nor2b_1
X_08343_ net335 VGND VPWR _00424_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[13\]
+ clknet_leaf_94_clk_regs sg13g2_dfrbpq_1
X_09037__945 VPWR VGND net1365 sg13g2_tiehi
X_05555_ _02238_ net3798 net1069 VPWR VGND sg13g2_nand2_1
X_08274_ net404 VGND VPWR _00355_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[8\]
+ clknet_leaf_101_clk_regs sg13g2_dfrbpq_1
X_07225_ net3600 net3587 net1086 _00950_ VPWR VGND sg13g2_mux2_1
X_05486_ _02184_ VPWR i_exotiny._1611_\[9\] VGND _02127_ _02183_ sg13g2_o21ai_1
X_08959__1023 VPWR VGND net1443 sg13g2_tiehi
X_07156_ net2198 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[13\]
+ net1008 _00904_ VPWR VGND sg13g2_mux2_1
XFILLER_106_748 VPWR VGND sg13g2_decap_8
XFILLER_105_214 VPWR VGND sg13g2_decap_8
X_06107_ net2756 _02523_ net958 _00280_ VPWR VGND sg13g2_mux2_1
X_07087_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[15\]
+ net3330 net915 _00842_ VPWR VGND sg13g2_mux2_1
X_06038_ net2766 net2562 net962 _00223_ VPWR VGND sg13g2_mux2_1
Xfanout1109 _01608_ net1109 VPWR VGND sg13g2_buf_8
XFILLER_102_965 VPWR VGND sg13g2_decap_8
XFILLER_101_464 VPWR VGND sg13g2_decap_8
XFILLER_74_315 VPWR VGND sg13g2_fill_2
XFILLER_59_367 VPWR VGND sg13g2_fill_1
X_07989_ net130 VGND VPWR net3444 i_exotiny._0369_\[14\] clknet_leaf_165_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_103_41 VPWR VGND sg13g2_fill_1
XFILLER_55_595 VPWR VGND sg13g2_decap_8
XFILLER_16_927 VPWR VGND sg13g2_fill_1
XFILLER_27_264 VPWR VGND sg13g2_fill_2
XFILLER_43_713 VPWR VGND sg13g2_decap_8
XFILLER_42_278 VPWR VGND sg13g2_fill_2
XFILLER_10_120 VPWR VGND sg13g2_fill_2
XFILLER_10_186 VPWR VGND sg13g2_fill_1
X_08779__1209 VPWR VGND net1629 sg13g2_tiehi
X_08815__1173 VPWR VGND net1593 sg13g2_tiehi
XFILLER_97_429 VPWR VGND sg13g2_decap_8
XFILLER_3_886 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_67_clk_regs clknet_5_24__leaf_clk_regs clknet_leaf_67_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_78_698 VPWR VGND sg13g2_fill_1
XFILLER_74_871 VPWR VGND sg13g2_fill_1
XFILLER_18_275 VPWR VGND sg13g2_fill_2
XFILLER_61_576 VPWR VGND sg13g2_fill_2
XFILLER_15_982 VPWR VGND sg13g2_decap_4
X_05340_ VGND VPWR _01832_ _01833_ _02064_ _02062_ sg13g2_a21oi_1
X_05271_ _01997_ _01792_ i_exotiny._0038_\[0\] _01785_ i_exotiny._0043_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_07010_ net3034 net3093 net921 _00777_ VPWR VGND sg13g2_mux2_1
XFILLER_45_0 VPWR VGND sg13g2_decap_4
XFILLER_102_217 VPWR VGND sg13g2_decap_8
X_08961_ net1441 VGND VPWR net2496 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[27\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
X_07912_ net736 VGND VPWR net2051 i_exotiny._1924_\[5\] clknet_leaf_33_clk_regs sg13g2_dfrbpq_1
X_08892_ net1510 VGND VPWR _00950_ i_exotiny.i_wb_spi.dat_rx_r\[22\] clknet_leaf_20_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_97_996 VPWR VGND sg13g2_decap_8
Xhold1815 i_exotiny.i_wdg_top.clk_div_inst.cnt\[8\] VPWR VGND net3642 sg13g2_dlygate4sd3_1
Xhold1804 _00678_ VPWR VGND net3631 sg13g2_dlygate4sd3_1
Xhold1826 _00010_ VPWR VGND net3653 sg13g2_dlygate4sd3_1
X_07843_ net3420 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[19\]
+ net983 _01316_ VPWR VGND sg13g2_mux2_1
Xhold1837 _00953_ VPWR VGND net3664 sg13g2_dlygate4sd3_1
Xhold1859 i_exotiny._1160_\[19\] VPWR VGND net3686 sg13g2_dlygate4sd3_1
Xhold1848 i_exotiny._0369_\[17\] VPWR VGND net3675 sg13g2_dlygate4sd3_1
X_07774_ net3321 net2132 net988 _01259_ VPWR VGND sg13g2_mux2_1
XFILLER_37_540 VPWR VGND sg13g2_fill_2
X_04986_ net1180 i_exotiny._6090_\[2\] i_exotiny._6090_\[3\] i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data[0]
+ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data[0]
+ _01706_ _01718_ VPWR VGND sg13g2_mux4_1
XFILLER_83_178 VPWR VGND sg13g2_fill_2
X_06725_ net3142 _02720_ _02757_ VPWR VGND sg13g2_nor2_1
X_06656_ _02696_ net2002 net1152 VPWR VGND sg13g2_nand2_1
X_05607_ net1116 i_exotiny._1924_\[2\] _02276_ VPWR VGND sg13g2_nor2b_1
X_06587_ net3509 net1153 _02648_ VPWR VGND sg13g2_nor2_1
XFILLER_21_930 VPWR VGND sg13g2_fill_2
X_08326_ net352 VGND VPWR _00407_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[28\]
+ clknet_leaf_83_clk_regs sg13g2_dfrbpq_1
X_08891__1091 VPWR VGND net1511 sg13g2_tiehi
XFILLER_20_451 VPWR VGND sg13g2_fill_1
X_05538_ VGND VPWR _01485_ _02220_ _02225_ _02224_ sg13g2_a21oi_1
X_08257_ net420 VGND VPWR _00338_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[24\]
+ clknet_leaf_49_clk_regs sg13g2_dfrbpq_1
X_05469_ _02168_ VPWR net31 VGND _02173_ _02174_ sg13g2_o21ai_1
X_08188_ net489 VGND VPWR _00269_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[19\]
+ clknet_leaf_70_clk_regs sg13g2_dfrbpq_1
X_07208_ VGND VPWR _01413_ net1088 _00939_ _02965_ sg13g2_a21oi_1
X_07139_ net1286 net1864 _00889_ VPWR VGND sg13g2_and2_1
XFILLER_106_545 VPWR VGND sg13g2_decap_8
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_58_23 VPWR VGND sg13g2_fill_2
XFILLER_59_153 VPWR VGND sg13g2_fill_1
XFILLER_58_78 VPWR VGND sg13g2_fill_1
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_101_261 VPWR VGND sg13g2_decap_8
XFILLER_48_838 VPWR VGND sg13g2_fill_2
XFILLER_90_605 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_185_clk_regs clknet_5_0__leaf_clk_regs clknet_leaf_185_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_15_223 VPWR VGND sg13g2_fill_2
XFILLER_71_874 VPWR VGND sg13g2_fill_2
XFILLER_15_245 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_114_clk_regs clknet_5_24__leaf_clk_regs clknet_leaf_114_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_8_923 VPWR VGND sg13g2_decap_8
XFILLER_12_974 VPWR VGND sg13g2_decap_8
XFILLER_97_204 VPWR VGND sg13g2_fill_2
X_08003__692 VPWR VGND net692 sg13g2_tiehi
X_09027__955 VPWR VGND net1375 sg13g2_tiehi
XFILLER_94_955 VPWR VGND sg13g2_decap_8
X_04840_ net3634 _01579_ _01580_ VPWR VGND sg13g2_nor2_2
X_04771_ _01522_ net3775 net1218 VPWR VGND sg13g2_nand2b_1
X_06510_ _02620_ net1142 net1160 _02621_ VPWR VGND sg13g2_a21o_2
XFILLER_0_63 VPWR VGND sg13g2_decap_4
X_07490_ net3555 net906 _03112_ VPWR VGND sg13g2_nor2_1
X_06441_ net2550 net2777 net937 _00528_ VPWR VGND sg13g2_mux2_1
X_06372_ net2522 net3135 net1030 _00502_ VPWR VGND sg13g2_mux2_1
X_08010__685 VPWR VGND net685 sg13g2_tiehi
X_09034__948 VPWR VGND net1368 sg13g2_tiehi
X_09160_ net822 VGND VPWR _01215_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[16\]
+ clknet_leaf_175_clk_regs sg13g2_dfrbpq_1
XFILLER_21_248 VPWR VGND sg13g2_fill_1
X_08111_ net583 VGND VPWR net2344 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[16\]
+ clknet_leaf_101_clk_regs sg13g2_dfrbpq_1
X_09091_ net1311 VGND VPWR net2707 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[11\]
+ clknet_leaf_145_clk_regs sg13g2_dfrbpq_1
X_05323_ _02045_ _02046_ _02047_ VPWR VGND sg13g2_nor2_1
X_08042_ net652 VGND VPWR net2904 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[11\]
+ clknet_leaf_56_clk_regs sg13g2_dfrbpq_1
X_05254_ _01980_ _01978_ _01979_ VPWR VGND sg13g2_nand2_1
Xhold912 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[11\]
+ VPWR VGND net2739 sg13g2_dlygate4sd3_1
Xhold901 _01192_ VPWR VGND net2728 sg13g2_dlygate4sd3_1
Xhold945 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[29\]
+ VPWR VGND net2772 sg13g2_dlygate4sd3_1
Xhold923 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[13\]
+ VPWR VGND net2750 sg13g2_dlygate4sd3_1
Xhold934 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[11\]
+ VPWR VGND net2761 sg13g2_dlygate4sd3_1
X_05185_ VGND VPWR _01913_ _01742_ _01736_ sg13g2_or2_1
XFILLER_89_727 VPWR VGND sg13g2_fill_1
Xhold989 _00081_ VPWR VGND net2816 sg13g2_dlygate4sd3_1
Xhold967 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[14\]
+ VPWR VGND net2794 sg13g2_dlygate4sd3_1
Xhold978 i_exotiny._0034_\[3\] VPWR VGND net2805 sg13g2_dlygate4sd3_1
Xhold956 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[10\]
+ VPWR VGND net2783 sg13g2_dlygate4sd3_1
X_08944_ net1458 VGND VPWR _01002_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[10\]
+ clknet_leaf_74_clk_regs sg13g2_dfrbpq_1
X_09080__902 VPWR VGND net1322 sg13g2_tiehi
Xhold1601 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[20\]
+ VPWR VGND net3428 sg13g2_dlygate4sd3_1
XFILLER_84_421 VPWR VGND sg13g2_fill_1
Xhold1612 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[17\]
+ VPWR VGND net3439 sg13g2_dlygate4sd3_1
Xhold1634 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[4\]
+ VPWR VGND net3461 sg13g2_dlygate4sd3_1
X_08875_ net1527 VGND VPWR _00933_ i_exotiny.i_wb_spi.dat_rx_r\[5\] clknet_leaf_26_clk_regs
+ sg13g2_dfrbpq_2
Xhold1623 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[14\]
+ VPWR VGND net3450 sg13g2_dlygate4sd3_1
XFILLER_28_37 VPWR VGND sg13g2_fill_1
Xhold1645 _01015_ VPWR VGND net3472 sg13g2_dlygate4sd3_1
XFILLER_84_443 VPWR VGND sg13g2_fill_1
Xhold1656 _00556_ VPWR VGND net3483 sg13g2_dlygate4sd3_1
XFILLER_72_605 VPWR VGND sg13g2_fill_2
XFILLER_56_134 VPWR VGND sg13g2_fill_2
Xhold1667 _00628_ VPWR VGND net3494 sg13g2_dlygate4sd3_1
Xhold1678 i_exotiny._0369_\[19\] VPWR VGND net3505 sg13g2_dlygate4sd3_1
X_07826_ net2162 i_exotiny._0022_\[2\] net984 _01299_ VPWR VGND sg13g2_mux2_1
X_07757_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[13\]
+ net2900 net991 _01242_ VPWR VGND sg13g2_mux2_1
Xhold1689 _00380_ VPWR VGND net3516 sg13g2_dlygate4sd3_1
XFILLER_85_999 VPWR VGND sg13g2_decap_8
XFILLER_38_871 VPWR VGND sg13g2_decap_4
X_04969_ _01695_ _01697_ _01693_ _01701_ VPWR VGND _01700_ sg13g2_nand4_1
X_06708_ net3719 net1102 _02743_ VPWR VGND sg13g2_nor2_1
XFILLER_53_863 VPWR VGND sg13g2_fill_1
X_07688_ net2176 net2974 net999 _01190_ VPWR VGND sg13g2_mux2_1
X_07901__47 VPWR VGND net47 sg13g2_tiehi
X_06639_ net1194 _02681_ _02682_ _00653_ VPWR VGND sg13g2_nor3_1
XFILLER_40_546 VPWR VGND sg13g2_fill_2
X_08309_ net369 VGND VPWR _00390_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[11\]
+ clknet_leaf_73_clk_regs sg13g2_dfrbpq_1
X_09289_ net1821 VGND VPWR _01344_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[15\]
+ clknet_leaf_168_clk_regs sg13g2_dfrbpq_1
XFILLER_106_342 VPWR VGND sg13g2_decap_8
XFILLER_5_959 VPWR VGND sg13g2_decap_8
XFILLER_69_33 VPWR VGND sg13g2_fill_1
XFILLER_62_126 VPWR VGND sg13g2_fill_1
XFILLER_90_479 VPWR VGND sg13g2_fill_1
XFILLER_31_502 VPWR VGND sg13g2_decap_8
XFILLER_43_384 VPWR VGND sg13g2_fill_1
XFILLER_15_1002 VPWR VGND sg13g2_fill_1
Xhold208 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[18\]
+ VPWR VGND net2035 sg13g2_dlygate4sd3_1
XFILLER_7_263 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_82_clk_regs clknet_5_27__leaf_clk_regs clknet_leaf_82_clk_regs VPWR VGND
+ sg13g2_buf_8
Xhold219 i_exotiny._1924_\[23\] VPWR VGND net2046 sg13g2_dlygate4sd3_1
XFILLER_98_502 VPWR VGND sg13g2_decap_8
XFILLER_4_981 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_11_clk_regs clknet_5_3__leaf_clk_regs clknet_leaf_11_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_100_507 VPWR VGND sg13g2_decap_8
X_06990_ net2803 net879 _02922_ _02926_ VPWR VGND sg13g2_mux2_1
X_05941_ net2168 net3295 net966 _00150_ VPWR VGND sg13g2_mux2_1
Xfanout1281 net1282 net1281 VPWR VGND sg13g2_buf_8
X_08660_ net1737 VGND VPWR _00728_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[29\]
+ clknet_leaf_148_clk_regs sg13g2_dfrbpq_1
X_05872_ VPWR VGND _01908_ _02458_ _02431_ _01496_ _02459_ _01911_ sg13g2_a221oi_1
XFILLER_39_657 VPWR VGND sg13g2_fill_2
Xfanout1270 net3754 net1270 VPWR VGND sg13g2_buf_8
X_04823_ net1866 net1854 net1864 _01562_ _01563_ VPWR VGND sg13g2_nor4_1
X_07611_ _03178_ net3649 _03176_ VPWR VGND sg13g2_xnor2_1
X_08591_ net1805 VGND VPWR _00663_ i_exotiny._6090_\[3\] clknet_leaf_9_clk_regs sg13g2_dfrbpq_2
X_07542_ VPWR _03134_ _03133_ VGND sg13g2_inv_1
X_04754_ net1174 _01454_ _01506_ VPWR VGND sg13g2_and2_1
XFILLER_61_170 VPWR VGND sg13g2_fill_1
X_04685_ net1281 VPWR _01444_ VGND _01364_ net3241 sg13g2_o21ai_1
X_07473_ net1211 net1239 _03008_ _01066_ VPWR VGND sg13g2_a21o_1
X_06424_ _02603_ net3611 net3689 VPWR VGND sg13g2_nand2_1
X_09212_ net767 VGND VPWR _01267_ i_exotiny._0023_\[2\] clknet_leaf_130_clk_regs sg13g2_dfrbpq_2
X_06355_ net2283 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[10\]
+ net1032 _00485_ VPWR VGND sg13g2_mux2_1
X_08774__1214 VPWR VGND net1634 sg13g2_tiehi
X_09143_ net839 VGND VPWR _01198_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[31\]
+ clknet_leaf_156_clk_regs sg13g2_dfrbpq_1
X_05306_ _02032_ _01630_ i_exotiny._0041_\[0\] _01615_ i_exotiny._0021_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_09074_ net1328 VGND VPWR _01129_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[14\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_06286_ net3332 net2963 net941 _00429_ VPWR VGND sg13g2_mux2_1
XFILLER_30_38 VPWR VGND sg13g2_fill_2
X_08025_ net669 VGND VPWR _00106_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[26\]
+ clknet_leaf_61_clk_regs sg13g2_dfrbpq_1
Xhold720 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[31\]
+ VPWR VGND net2547 sg13g2_dlygate4sd3_1
X_05237_ _01958_ _01959_ _01957_ _01965_ VPWR VGND _01964_ sg13g2_nand4_1
Xhold764 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[27\]
+ VPWR VGND net2591 sg13g2_dlygate4sd3_1
Xhold731 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[19\]
+ VPWR VGND net2558 sg13g2_dlygate4sd3_1
Xhold753 _01212_ VPWR VGND net2580 sg13g2_dlygate4sd3_1
Xhold742 _01214_ VPWR VGND net2569 sg13g2_dlygate4sd3_1
XFILLER_2_929 VPWR VGND sg13g2_decap_8
X_05168_ VPWR VGND _01870_ net1110 _01845_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[2\]
+ _01898_ net1107 sg13g2_a221oi_1
XFILLER_104_846 VPWR VGND sg13g2_decap_8
XFILLER_89_524 VPWR VGND sg13g2_fill_2
Xhold775 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[15\]
+ VPWR VGND net2602 sg13g2_dlygate4sd3_1
Xhold786 i_exotiny._0027_\[2\] VPWR VGND net2613 sg13g2_dlygate4sd3_1
XFILLER_1_428 VPWR VGND sg13g2_fill_2
Xhold797 _00607_ VPWR VGND net2624 sg13g2_dlygate4sd3_1
XFILLER_103_367 VPWR VGND sg13g2_decap_8
XFILLER_77_719 VPWR VGND sg13g2_fill_1
X_05099_ net1248 _01823_ _01829_ VPWR VGND sg13g2_and2_1
X_08927_ net1475 VGND VPWR _00985_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[25\]
+ clknet_leaf_113_clk_regs sg13g2_dfrbpq_1
X_08549__107 VPWR VGND net107 sg13g2_tiehi
Xhold1442 i_exotiny._0028_\[0\] VPWR VGND net3269 sg13g2_dlygate4sd3_1
Xhold1420 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[7\]
+ VPWR VGND net3247 sg13g2_dlygate4sd3_1
X_08858_ net1548 VGND VPWR _00916_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[25\]
+ clknet_leaf_186_clk_regs sg13g2_dfrbpq_1
Xhold1431 _00457_ VPWR VGND net3258 sg13g2_dlygate4sd3_1
XFILLER_85_785 VPWR VGND sg13g2_fill_2
Xhold1453 _00267_ VPWR VGND net3280 sg13g2_dlygate4sd3_1
Xhold1464 i_exotiny._0039_\[2\] VPWR VGND net3291 sg13g2_dlygate4sd3_1
Xhold1486 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[22\]
+ VPWR VGND net3313 sg13g2_dlygate4sd3_1
Xhold1475 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[28\]
+ VPWR VGND net3302 sg13g2_dlygate4sd3_1
X_07809_ net2345 net2781 net891 _01288_ VPWR VGND sg13g2_mux2_1
Xhold1497 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[28\]
+ VPWR VGND net3324 sg13g2_dlygate4sd3_1
X_08789_ net1619 VGND VPWR net3414 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[20\]
+ clknet_leaf_167_clk_regs sg13g2_dfrbpq_1
XFILLER_44_115 VPWR VGND sg13g2_fill_1
XFILLER_41_877 VPWR VGND sg13g2_fill_1
X_09017__965 VPWR VGND net1385 sg13g2_tiehi
XFILLER_41_899 VPWR VGND sg13g2_fill_1
X_08000__695 VPWR VGND net695 sg13g2_tiehi
XFILLER_76_763 VPWR VGND sg13g2_fill_2
X_09024__958 VPWR VGND net1378 sg13g2_tiehi
XFILLER_75_251 VPWR VGND sg13g2_fill_1
Xhold80 i_exotiny._1924_\[4\] VPWR VGND net1907 sg13g2_dlygate4sd3_1
XFILLER_63_402 VPWR VGND sg13g2_fill_2
Xhold91 i_exotiny._1924_\[28\] VPWR VGND net1918 sg13g2_dlygate4sd3_1
XFILLER_64_947 VPWR VGND sg13g2_fill_1
XFILLER_63_446 VPWR VGND sg13g2_fill_2
XFILLER_91_1015 VPWR VGND sg13g2_decap_8
XFILLER_43_192 VPWR VGND sg13g2_fill_2
X_09070__912 VPWR VGND net1332 sg13g2_tiehi
X_06140_ net2658 net2333 net1046 _00309_ VPWR VGND sg13g2_mux2_1
X_06071_ VGND VPWR _02518_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[4\]
+ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.rd_i\[3\] sg13g2_or2_1
XFILLER_99_811 VPWR VGND sg13g2_fill_1
XFILLER_6_84 VPWR VGND sg13g2_fill_2
X_05022_ _01754_ i_exotiny._0079_\[2\] i_exotiny._0079_\[3\] VPWR VGND sg13g2_nand2_2
XFILLER_99_877 VPWR VGND sg13g2_decap_8
XFILLER_100_304 VPWR VGND sg13g2_decap_8
XFILLER_98_376 VPWR VGND sg13g2_decap_8
X_06973_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[15\]
+ net2280 net1020 _00746_ VPWR VGND sg13g2_mux2_1
XFILLER_6_1011 VPWR VGND sg13g2_decap_8
X_05924_ net3120 _02480_ net975 _00140_ VPWR VGND sg13g2_mux2_1
X_08712_ net1696 VGND VPWR _00770_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[7\]
+ clknet_leaf_117_clk_regs sg13g2_dfrbpq_1
X_08828__1160 VPWR VGND net1580 sg13g2_tiehi
XFILLER_66_251 VPWR VGND sg13g2_fill_2
XFILLER_66_240 VPWR VGND sg13g2_fill_2
XFILLER_55_914 VPWR VGND sg13g2_fill_1
XFILLER_82_722 VPWR VGND sg13g2_fill_2
X_08643_ net1754 VGND VPWR net3381 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[12\]
+ clknet_leaf_146_clk_regs sg13g2_dfrbpq_1
X_05855_ _02438_ VPWR _02444_ VGND _02442_ _02443_ sg13g2_o21ai_1
X_05786_ _02408_ i_exotiny._2034_\[9\] _00026_ VPWR VGND sg13g2_nand2_1
XFILLER_70_906 VPWR VGND sg13g2_fill_1
X_04806_ net3789 net1234 _01465_ i_exotiny._2160_ VGND VPWR _01551_ sg13g2_nor4_2
X_08574_ net56 VGND VPWR net3156 i_exotiny._0314_\[19\] clknet_leaf_179_clk_regs sg13g2_dfrbpq_1
XFILLER_82_799 VPWR VGND sg13g2_fill_2
X_04737_ VGND VPWR _01493_ _01486_ i_exotiny.i_wb_qspi_mem.cnt_r\[2\] sg13g2_or2_1
X_07525_ _03119_ VPWR _01100_ VGND _03120_ _03121_ sg13g2_o21ai_1
XFILLER_50_641 VPWR VGND sg13g2_fill_1
XFILLER_23_899 VPWR VGND sg13g2_fill_1
X_07456_ _03093_ VPWR _01059_ VGND net1080 _03092_ sg13g2_o21ai_1
X_08479__201 VPWR VGND net201 sg13g2_tiehi
X_04668_ net1249 net1247 net1243 _01429_ VPWR VGND sg13g2_nor3_2
X_04599_ net3567 _01361_ VPWR VGND sg13g2_inv_4
X_07387_ i_exotiny._0369_\[30\] net1214 _03041_ VPWR VGND sg13g2_and2_1
X_06407_ _02590_ net2014 net1071 VPWR VGND sg13g2_nand2_1
X_06338_ i_exotiny._0014_\[2\] net877 _02558_ _02562_ VPWR VGND sg13g2_mux2_1
X_09126_ net856 VGND VPWR net3182 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[14\]
+ clknet_leaf_156_clk_regs sg13g2_dfrbpq_1
XFILLER_41_59 VPWR VGND sg13g2_fill_1
X_06269_ net2119 i_exotiny._0016_\[1\] net939 _00412_ VPWR VGND sg13g2_mux2_1
X_09057_ net1345 VGND VPWR _01112_ i_exotiny._1652_\[0\] clknet_leaf_22_clk_regs sg13g2_dfrbpq_1
X_08008_ net687 VGND VPWR _00089_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[9\]
+ clknet_leaf_66_clk_regs sg13g2_dfrbpq_1
XFILLER_104_621 VPWR VGND sg13g2_decap_8
Xhold572 _00989_ VPWR VGND net2399 sg13g2_dlygate4sd3_1
Xhold550 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[14\]
+ VPWR VGND net2377 sg13g2_dlygate4sd3_1
Xhold561 _01222_ VPWR VGND net2388 sg13g2_dlygate4sd3_1
Xhold583 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[4\]
+ VPWR VGND net2410 sg13g2_dlygate4sd3_1
XFILLER_104_643 VPWR VGND sg13g2_decap_8
Xhold594 _01179_ VPWR VGND net2421 sg13g2_dlygate4sd3_1
XFILLER_103_164 VPWR VGND sg13g2_decap_8
XFILLER_89_398 VPWR VGND sg13g2_fill_1
XFILLER_100_882 VPWR VGND sg13g2_decap_8
Xhold1261 _00385_ VPWR VGND net3088 sg13g2_dlygate4sd3_1
Xhold1250 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[30\]
+ VPWR VGND net3077 sg13g2_dlygate4sd3_1
Xhold1283 _00802_ VPWR VGND net3110 sg13g2_dlygate4sd3_1
Xhold1294 _00140_ VPWR VGND net3121 sg13g2_dlygate4sd3_1
Xhold1272 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[12\]
+ VPWR VGND net3099 sg13g2_dlygate4sd3_1
XFILLER_17_159 VPWR VGND sg13g2_fill_2
XFILLER_45_468 VPWR VGND sg13g2_fill_1
XFILLER_14_833 VPWR VGND sg13g2_fill_1
XFILLER_25_181 VPWR VGND sg13g2_fill_2
XFILLER_41_630 VPWR VGND sg13g2_fill_2
XFILLER_12_1016 VPWR VGND sg13g2_decap_8
XFILLER_12_1027 VPWR VGND sg13g2_fill_2
X_08139__546 VPWR VGND net546 sg13g2_tiehi
XFILLER_68_527 VPWR VGND sg13g2_fill_1
XFILLER_96_858 VPWR VGND sg13g2_decap_8
XFILLER_95_335 VPWR VGND sg13g2_decap_8
XFILLER_83_508 VPWR VGND sg13g2_fill_1
XFILLER_48_240 VPWR VGND sg13g2_fill_1
XFILLER_91_552 VPWR VGND sg13g2_fill_1
X_05640_ net1124 i_exotiny._1924_\[10\] _02301_ VPWR VGND sg13g2_nor2b_1
X_05571_ net1234 i_exotiny._0327_\[0\] _02251_ VPWR VGND sg13g2_xor2_1
X_07310_ net2495 _02983_ net911 _01023_ VPWR VGND sg13g2_mux2_1
X_08290_ net388 VGND VPWR net2480 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[24\]
+ clknet_leaf_99_clk_regs sg13g2_dfrbpq_1
X_08146__539 VPWR VGND net539 sg13g2_tiehi
X_07241_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[8\]
+ net3314 net1007 _00964_ VPWR VGND sg13g2_mux2_1
Xclkbuf_4_0_0_clk_regs clknet_0_clk_regs clknet_4_0_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_75_0 VPWR VGND sg13g2_fill_1
X_07172_ _02949_ net3533 net1011 _00919_ VPWR VGND sg13g2_mux2_1
XFILLER_9_892 VPWR VGND sg13g2_fill_1
X_06123_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[14\]
+ net2691 net1045 _00292_ VPWR VGND sg13g2_mux2_1
X_08122__572 VPWR VGND net572 sg13g2_tiehi
X_06054_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[26\]
+ net2699 net961 _00239_ VPWR VGND sg13g2_mux2_1
X_05005_ _01708_ _01734_ _01391_ _01737_ VPWR VGND _01735_ sg13g2_nand4_1
X_06956_ _02492_ _02518_ _02922_ VPWR VGND sg13g2_nor2_2
X_09007__975 VPWR VGND net1395 sg13g2_tiehi
XFILLER_95_891 VPWR VGND sg13g2_decap_8
X_05907_ net2931 net3392 net975 _00124_ VPWR VGND sg13g2_mux2_1
X_06887_ net3387 net1189 _02893_ VPWR VGND sg13g2_nor2_1
X_08626_ net741 VGND VPWR net2572 i_exotiny.core_res_en_n clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_2
X_05838_ VGND VPWR net1243 _01605_ _02427_ _01816_ sg13g2_a21oi_1
X_05769_ _02397_ net1126 net2033 net1144 net3528 VPWR VGND sg13g2_a22oi_1
X_08557_ net98 VGND VPWR net3408 i_exotiny._0314_\[2\] clknet_leaf_13_clk_regs sg13g2_dfrbpq_2
X_08488_ net192 VGND VPWR _00562_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[8\]
+ clknet_leaf_108_clk_regs sg13g2_dfrbpq_1
X_07508_ net3220 net3318 net902 _01091_ VPWR VGND sg13g2_mux2_1
XFILLER_7_807 VPWR VGND sg13g2_fill_1
X_07439_ VGND VPWR net3558 net1082 _03082_ _03077_ sg13g2_a21oi_1
X_08851__1135 VPWR VGND net1555 sg13g2_tiehi
X_09109_ net1293 VGND VPWR _01164_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[29\]
+ clknet_leaf_153_clk_regs sg13g2_dfrbpq_1
X_09014__968 VPWR VGND net1388 sg13g2_tiehi
XFILLER_105_930 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_139_clk_regs clknet_5_17__leaf_clk_regs clknet_leaf_139_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_2_512 VPWR VGND sg13g2_fill_1
XFILLER_2_523 VPWR VGND sg13g2_fill_2
X_07997__532 VPWR VGND net532 sg13g2_tiehi
Xhold380 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[6\]
+ VPWR VGND net2207 sg13g2_dlygate4sd3_1
Xhold391 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[13\]
+ VPWR VGND net2218 sg13g2_dlygate4sd3_1
XFILLER_104_495 VPWR VGND sg13g2_decap_8
X_09060__922 VPWR VGND net1342 sg13g2_tiehi
XFILLER_92_305 VPWR VGND sg13g2_decap_8
Xfanout893 net895 net893 VPWR VGND sg13g2_buf_8
Xfanout882 net884 net882 VPWR VGND sg13g2_buf_8
XFILLER_46_700 VPWR VGND sg13g2_decap_8
Xhold1080 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[14\]
+ VPWR VGND net2907 sg13g2_dlygate4sd3_1
X_08595__1381 VPWR VGND net1801 sg13g2_tiehi
Xhold1091 _01138_ VPWR VGND net2918 sg13g2_dlygate4sd3_1
XFILLER_60_246 VPWR VGND sg13g2_fill_1
XFILLER_33_449 VPWR VGND sg13g2_fill_2
X_09169__813 VPWR VGND net813 sg13g2_tiehi
XFILLER_95_121 VPWR VGND sg13g2_fill_2
X_06810_ net1171 VPWR _02829_ VGND net1937 net1185 sg13g2_o21ai_1
X_07790_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[4\]
+ net2071 net893 _01269_ VPWR VGND sg13g2_mux2_1
X_08469__211 VPWR VGND net211 sg13g2_tiehi
XFILLER_97_1010 VPWR VGND sg13g2_decap_8
X_09176__806 VPWR VGND net806 sg13g2_tiehi
X_06741_ VGND VPWR net2331 net1130 _02771_ _02770_ sg13g2_a21oi_1
XFILLER_37_711 VPWR VGND sg13g2_fill_2
XFILLER_92_861 VPWR VGND sg13g2_fill_2
XFILLER_36_232 VPWR VGND sg13g2_fill_2
X_08411_ net274 VGND VPWR net2284 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[10\]
+ clknet_leaf_97_clk_regs sg13g2_dfrbpq_1
X_06672_ _02710_ _02707_ _02709_ VPWR VGND sg13g2_nand2b_1
X_05623_ net1895 net1065 _02288_ VPWR VGND sg13g2_nor2_1
X_08342_ net336 VGND VPWR net2508 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[12\]
+ clknet_leaf_96_clk_regs sg13g2_dfrbpq_1
X_05554_ _02235_ VPWR i_exotiny._1611_\[29\] VGND _02219_ _02237_ sg13g2_o21ai_1
X_08273_ net405 VGND VPWR net3496 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[7\]
+ clknet_leaf_99_clk_regs sg13g2_dfrbpq_1
X_05485_ _02184_ net3601 net1071 VPWR VGND sg13g2_nand2_1
X_08632__1345 VPWR VGND net1765 sg13g2_tiehi
X_07224_ net3644 net3600 net1086 _00949_ VPWR VGND sg13g2_mux2_1
X_08476__204 VPWR VGND net204 sg13g2_tiehi
X_07155_ net2323 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[12\]
+ net1011 _00903_ VPWR VGND sg13g2_mux2_1
XFILLER_106_727 VPWR VGND sg13g2_decap_8
X_06106_ i_exotiny._0038_\[2\] net878 _02519_ _02523_ VPWR VGND sg13g2_mux2_1
X_07086_ net3364 net3367 net917 _00841_ VPWR VGND sg13g2_mux2_1
X_06037_ net3500 net3485 net962 _00222_ VPWR VGND sg13g2_mux2_1
X_08196__481 VPWR VGND net481 sg13g2_tiehi
XFILLER_102_944 VPWR VGND sg13g2_decap_8
XFILLER_99_493 VPWR VGND sg13g2_decap_8
X_09044__939 VPWR VGND net1359 sg13g2_tiehi
XFILLER_101_443 VPWR VGND sg13g2_decap_8
X_07988_ net129 VGND VPWR net2998 i_exotiny._0369_\[13\] clknet_leaf_14_clk_regs sg13g2_dfrbpq_2
X_06939_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[19\]
+ net2315 net927 _00718_ VPWR VGND sg13g2_mux2_1
XFILLER_42_202 VPWR VGND sg13g2_fill_2
X_08609_ net1787 VGND VPWR _00681_ i_exotiny._1617_\[1\] clknet_leaf_22_clk_regs sg13g2_dfrbpq_2
XFILLER_42_246 VPWR VGND sg13g2_fill_1
X_08583__1396 VPWR VGND net1816 sg13g2_tiehi
XFILLER_98_909 VPWR VGND sg13g2_decap_8
XFILLER_97_408 VPWR VGND sg13g2_decap_8
XFILLER_3_865 VPWR VGND sg13g2_decap_8
X_08787__1201 VPWR VGND net1621 sg13g2_tiehi
XFILLER_104_292 VPWR VGND sg13g2_decap_8
XFILLER_66_817 VPWR VGND sg13g2_fill_1
X_08136__549 VPWR VGND net549 sg13g2_tiehi
X_08710__1278 VPWR VGND net1698 sg13g2_tiehi
Xclkbuf_leaf_36_clk_regs clknet_5_11__leaf_clk_regs clknet_leaf_36_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_19_799 VPWR VGND sg13g2_fill_1
XFILLER_33_202 VPWR VGND sg13g2_fill_2
XFILLER_37_91 VPWR VGND sg13g2_fill_2
X_08112__582 VPWR VGND net582 sg13g2_tiehi
XFILLER_18_1000 VPWR VGND sg13g2_fill_2
XFILLER_105_1014 VPWR VGND sg13g2_decap_8
XFILLER_30_997 VPWR VGND sg13g2_fill_2
X_05270_ _01993_ _01994_ _01991_ _01996_ VPWR VGND _01995_ sg13g2_nand4_1
XFILLER_89_909 VPWR VGND sg13g2_fill_1
X_08960_ net1442 VGND VPWR net2291 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[26\]
+ clknet_leaf_74_clk_regs sg13g2_dfrbpq_1
XFILLER_96_430 VPWR VGND sg13g2_decap_8
X_07911_ net737 VGND VPWR net1908 i_exotiny._1924_\[4\] clknet_leaf_33_clk_regs sg13g2_dfrbpq_1
X_08891_ net1511 VGND VPWR _00949_ i_exotiny.i_wb_spi.dat_rx_r\[21\] clknet_leaf_63_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_38_0 VPWR VGND sg13g2_fill_1
XFILLER_97_975 VPWR VGND sg13g2_decap_8
XFILLER_96_452 VPWR VGND sg13g2_fill_2
Xhold1827 i_exotiny.i_wb_spi.dat_rx_r\[4\] VPWR VGND net3654 sg13g2_dlygate4sd3_1
Xhold1805 i_exotiny._6090_\[0\] VPWR VGND net3632 sg13g2_dlygate4sd3_1
Xhold1816 i_exotiny._0369_\[14\] VPWR VGND net3643 sg13g2_dlygate4sd3_1
X_07842_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[22\]
+ net2922 net984 _01315_ VPWR VGND sg13g2_mux2_1
Xhold1838 i_exotiny._0315_\[12\] VPWR VGND net3665 sg13g2_dlygate4sd3_1
Xhold1849 i_exotiny._1611_\[13\] VPWR VGND net3676 sg13g2_dlygate4sd3_1
X_07773_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[29\]
+ net2696 net991 _01258_ VPWR VGND sg13g2_mux2_1
XFILLER_65_850 VPWR VGND sg13g2_fill_2
X_04985_ VGND VPWR net1250 i_exotiny._0550_ _01717_ _01716_ sg13g2_a21oi_1
XFILLER_65_883 VPWR VGND sg13g2_fill_2
XFILLER_65_872 VPWR VGND sg13g2_fill_1
X_06724_ _02756_ VPWR _00664_ VGND net1137 _02755_ sg13g2_o21ai_1
XFILLER_52_511 VPWR VGND sg13g2_fill_2
X_09004__978 VPWR VGND net1398 sg13g2_tiehi
XFILLER_80_831 VPWR VGND sg13g2_fill_1
X_09287__1405 VPWR VGND net1825 sg13g2_tiehi
X_06655_ VGND VPWR _02687_ _02695_ _00656_ net1195 sg13g2_a21oi_1
XFILLER_24_235 VPWR VGND sg13g2_fill_1
XFILLER_80_864 VPWR VGND sg13g2_fill_1
X_05606_ VGND VPWR net1060 _02275_ _00027_ _02274_ sg13g2_a21oi_1
XFILLER_24_257 VPWR VGND sg13g2_fill_2
X_08325_ net353 VGND VPWR _00406_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[27\]
+ clknet_leaf_73_clk_regs sg13g2_dfrbpq_1
X_06586_ net3476 net1159 _02647_ VPWR VGND sg13g2_nor2_1
XFILLER_33_780 VPWR VGND sg13g2_fill_1
X_05537_ VPWR VGND _02223_ _02221_ _02222_ _01484_ _02224_ _01513_ sg13g2_a221oi_1
X_09050__932 VPWR VGND net1352 sg13g2_tiehi
X_08256_ net421 VGND VPWR _00337_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[23\]
+ clknet_leaf_57_clk_regs sg13g2_dfrbpq_1
X_05468_ net1264 VPWR _02174_ VGND i_exotiny._1619_\[3\] _02138_ sg13g2_o21ai_1
Xclkbuf_5_19__f_clk_regs clknet_4_9_0_clk_regs clknet_5_19__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08187_ net490 VGND VPWR net2414 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[18\]
+ clknet_leaf_68_clk_regs sg13g2_dfrbpq_1
X_07207_ net2105 net1088 _02965_ VPWR VGND sg13g2_nor2_1
X_08908__1074 VPWR VGND net1494 sg13g2_tiehi
XFILLER_106_524 VPWR VGND sg13g2_decap_8
X_07138_ net1286 net1844 _00888_ VPWR VGND sg13g2_and2_1
X_05399_ net1113 _02113_ _02114_ i_exotiny._2043_\[3\] VPWR VGND sg13g2_nor3_1
X_09228__751 VPWR VGND net751 sg13g2_tiehi
X_07069_ _02939_ net3047 net1014 _00826_ VPWR VGND sg13g2_mux2_1
XFILLER_99_290 VPWR VGND sg13g2_decap_8
XFILLER_102_752 VPWR VGND sg13g2_decap_8
XFILLER_101_240 VPWR VGND sg13g2_decap_8
XFILLER_88_986 VPWR VGND sg13g2_decap_8
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_74_157 VPWR VGND sg13g2_fill_1
X_09159__823 VPWR VGND net823 sg13g2_tiehi
XFILLER_83_680 VPWR VGND sg13g2_fill_1
XFILLER_16_736 VPWR VGND sg13g2_fill_2
XFILLER_71_886 VPWR VGND sg13g2_fill_2
XFILLER_15_268 VPWR VGND sg13g2_fill_1
X_09235__744 VPWR VGND net744 sg13g2_tiehi
XFILLER_12_953 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_154_clk_regs clknet_5_18__leaf_clk_regs clknet_leaf_154_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08459__221 VPWR VGND net221 sg13g2_tiehi
XFILLER_8_979 VPWR VGND sg13g2_decap_8
XFILLER_87_1020 VPWR VGND sg13g2_decap_8
X_09166__816 VPWR VGND net816 sg13g2_tiehi
XFILLER_48_1026 VPWR VGND sg13g2_fill_2
XFILLER_3_662 VPWR VGND sg13g2_fill_1
XFILLER_31_7 VPWR VGND sg13g2_decap_4
XFILLER_94_934 VPWR VGND sg13g2_decap_8
XFILLER_66_636 VPWR VGND sg13g2_fill_1
XFILLER_66_614 VPWR VGND sg13g2_fill_2
XFILLER_38_316 VPWR VGND sg13g2_fill_2
X_08466__214 VPWR VGND net214 sg13g2_tiehi
XFILLER_81_617 VPWR VGND sg13g2_fill_1
X_04770_ _01521_ net3830 _01519_ VPWR VGND sg13g2_nand2_2
XFILLER_0_42 VPWR VGND sg13g2_decap_8
X_09173__809 VPWR VGND net809 sg13g2_tiehi
X_06440_ net2232 net3037 net934 _00527_ VPWR VGND sg13g2_mux2_1
X_08186__491 VPWR VGND net491 sg13g2_tiehi
X_06371_ net2718 net2196 net1031 _00501_ VPWR VGND sg13g2_mux2_1
X_09090_ net1312 VGND VPWR net2687 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[10\]
+ clknet_leaf_142_clk_regs sg13g2_dfrbpq_1
XFILLER_30_772 VPWR VGND sg13g2_fill_2
X_05322_ _01831_ _02043_ _02044_ _02046_ VPWR VGND sg13g2_nor3_1
X_08110_ net584 VGND VPWR _00191_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[15\]
+ clknet_leaf_125_clk_regs sg13g2_dfrbpq_1
X_08041_ net653 VGND VPWR net2818 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[10\]
+ clknet_leaf_52_clk_regs sg13g2_dfrbpq_1
X_05253_ _01977_ _01976_ _01972_ _01979_ VPWR VGND sg13g2_a21o_2
Xhold902 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[26\]
+ VPWR VGND net2729 sg13g2_dlygate4sd3_1
Xhold913 _00325_ VPWR VGND net2740 sg13g2_dlygate4sd3_1
X_08473__207 VPWR VGND net207 sg13g2_tiehi
Xhold946 _00173_ VPWR VGND net2773 sg13g2_dlygate4sd3_1
X_08868__1116 VPWR VGND net1536 sg13g2_tiehi
Xhold935 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[8\]
+ VPWR VGND net2762 sg13g2_dlygate4sd3_1
Xhold924 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[14\]
+ VPWR VGND net2751 sg13g2_dlygate4sd3_1
X_05184_ _01912_ _01908_ _01910_ _01835_ _01834_ VPWR VGND sg13g2_a22oi_1
Xhold979 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[29\]
+ VPWR VGND net2806 sg13g2_dlygate4sd3_1
Xhold957 _00709_ VPWR VGND net2784 sg13g2_dlygate4sd3_1
Xhold968 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[29\]
+ VPWR VGND net2795 sg13g2_dlygate4sd3_1
X_08943_ net1459 VGND VPWR net2068 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[9\]
+ clknet_leaf_74_clk_regs sg13g2_dfrbpq_1
XFILLER_97_772 VPWR VGND sg13g2_fill_2
X_08193__484 VPWR VGND net484 sg13g2_tiehi
X_08874_ net1528 VGND VPWR net3557 i_exotiny.i_wb_spi.dat_rx_r\[4\] clknet_leaf_27_clk_regs
+ sg13g2_dfrbpq_1
Xhold1602 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[4\]
+ VPWR VGND net3429 sg13g2_dlygate4sd3_1
Xhold1624 _00296_ VPWR VGND net3451 sg13g2_dlygate4sd3_1
Xhold1613 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[22\]
+ VPWR VGND net3440 sg13g2_dlygate4sd3_1
Xhold1635 i_exotiny._0314_\[14\] VPWR VGND net3462 sg13g2_dlygate4sd3_1
XFILLER_85_978 VPWR VGND sg13g2_decap_8
Xhold1668 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[7\]
+ VPWR VGND net3495 sg13g2_dlygate4sd3_1
Xhold1646 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[16\]
+ VPWR VGND net3473 sg13g2_dlygate4sd3_1
X_07825_ net3491 i_exotiny._0022_\[1\] net985 _01298_ VPWR VGND sg13g2_mux2_1
Xhold1657 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[8\]
+ VPWR VGND net3484 sg13g2_dlygate4sd3_1
X_07756_ net2404 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[8\]
+ net991 _01241_ VPWR VGND sg13g2_mux2_1
Xhold1679 i_exotiny._1611_\[15\] VPWR VGND net3506 sg13g2_dlygate4sd3_1
X_04968_ VGND VPWR i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[2\] _01696_ _01700_
+ _01699_ sg13g2_a21oi_1
X_07898__44 VPWR VGND net44 sg13g2_tiehi
X_06707_ i_exotiny._0369_\[2\] net3574 net1193 _02742_ VPWR VGND sg13g2_mux2_1
X_04899_ net1222 _01617_ _01623_ _01631_ VPWR VGND sg13g2_nor3_2
XFILLER_25_577 VPWR VGND sg13g2_fill_1
X_07687_ net2499 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[26\]
+ net1001 _01189_ VPWR VGND sg13g2_mux2_1
XFILLER_13_728 VPWR VGND sg13g2_fill_2
X_06638_ net2002 net1153 _02682_ VPWR VGND sg13g2_nor2_1
X_06569_ net3407 net1155 _02636_ VPWR VGND sg13g2_nor2_1
X_08308_ net370 VGND VPWR _00389_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[10\]
+ clknet_leaf_72_clk_regs sg13g2_dfrbpq_1
X_09288_ net1823 VGND VPWR net3251 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[14\]
+ clknet_leaf_171_clk_regs sg13g2_dfrbpq_1
X_08239_ net438 VGND VPWR _00320_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[6\]
+ clknet_leaf_48_clk_regs sg13g2_dfrbpq_1
XFILLER_5_938 VPWR VGND sg13g2_decap_8
XFILLER_106_321 VPWR VGND sg13g2_decap_8
Xclkbuf_4_13_0_clk_regs clknet_0_clk_regs clknet_4_13_0_clk_regs VPWR VGND sg13g2_buf_8
XFILLER_106_398 VPWR VGND sg13g2_decap_8
X_08102__592 VPWR VGND net592 sg13g2_tiehi
XFILLER_91_959 VPWR VGND sg13g2_decap_8
XFILLER_16_599 VPWR VGND sg13g2_fill_1
XFILLER_43_374 VPWR VGND sg13g2_fill_2
XFILLER_102_1028 VPWR VGND sg13g2_fill_1
XFILLER_8_776 VPWR VGND sg13g2_fill_1
Xhold209 _01006_ VPWR VGND net2036 sg13g2_dlygate4sd3_1
XFILLER_4_960 VPWR VGND sg13g2_decap_8
XFILLER_98_525 VPWR VGND sg13g2_fill_1
X_08864__1122 VPWR VGND net1542 sg13g2_tiehi
Xclkbuf_leaf_51_clk_regs clknet_5_15__leaf_clk_regs clknet_leaf_51_clk_regs VPWR VGND
+ sg13g2_buf_8
X_05940_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[5\]
+ net2418 net969 _00149_ VPWR VGND sg13g2_mux2_1
XFILLER_94_764 VPWR VGND sg13g2_fill_1
Xfanout1282 net1291 net1282 VPWR VGND sg13g2_buf_8
Xfanout1271 net1274 net1271 VPWR VGND sg13g2_buf_8
X_05871_ _01498_ _01910_ _02458_ VPWR VGND sg13g2_nor2_1
Xfanout1260 net1261 net1260 VPWR VGND sg13g2_buf_8
X_04822_ i_exotiny.i_wb_spi.state_r\[24\] i_exotiny.i_wb_spi.state_r\[27\] i_exotiny.i_wb_spi.state_r\[26\]
+ i_exotiny.i_wb_spi.state_r\[29\] _01562_ VPWR VGND sg13g2_or4_1
X_07610_ _03176_ net3723 _01129_ VPWR VGND sg13g2_nor2_1
X_09040__942 VPWR VGND net1362 sg13g2_tiehi
X_08590_ net1806 VGND VPWR net3720 i_exotiny._6090_\[2\] clknet_leaf_8_clk_regs sg13g2_dfrbpq_2
XFILLER_93_296 VPWR VGND sg13g2_decap_8
X_07541_ _03133_ net3466 net1290 VPWR VGND sg13g2_nand2_2
X_04753_ _01488_ net3651 net1226 _00006_ VPWR VGND sg13g2_a21o_1
X_09218__761 VPWR VGND net761 sg13g2_tiehi
X_04684_ i_exotiny._1265_ _01443_ VPWR VGND sg13g2_inv_2
X_07472_ net1211 net1241 _03044_ _01065_ VPWR VGND sg13g2_a21o_1
X_06423_ VGND VPWR net3430 _02595_ _02602_ net1227 sg13g2_a21oi_1
X_09211_ net768 VGND VPWR net3204 i_exotiny._0023_\[1\] clknet_leaf_128_clk_regs sg13g2_dfrbpq_2
X_06354_ net3354 net3379 net1028 _00484_ VPWR VGND sg13g2_mux2_1
X_09142_ net840 VGND VPWR _01197_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[30\]
+ clknet_leaf_157_clk_regs sg13g2_dfrbpq_1
X_05305_ _02031_ _01648_ i_exotiny._0033_\[0\] _01637_ i_exotiny._0024_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_09073_ net1329 VGND VPWR net3237 i_exotiny.i_wdg_top.clk_div_inst.cnt\[13\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_06285_ net2367 net2797 net940 _00428_ VPWR VGND sg13g2_mux2_1
Xhold721 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[8\]
+ VPWR VGND net2548 sg13g2_dlygate4sd3_1
X_08024_ net670 VGND VPWR _00105_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[25\]
+ clknet_leaf_67_clk_regs sg13g2_dfrbpq_1
X_05236_ _01960_ _01961_ _01962_ _01963_ _01964_ VPWR VGND sg13g2_and4_1
X_09149__833 VPWR VGND net833 sg13g2_tiehi
Xhold710 _01320_ VPWR VGND net2537 sg13g2_dlygate4sd3_1
Xhold754 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[18\]
+ VPWR VGND net2581 sg13g2_dlygate4sd3_1
Xhold732 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[27\]
+ VPWR VGND net2559 sg13g2_dlygate4sd3_1
Xhold743 i_exotiny.i_rstctl.wdg_res_n VPWR VGND net2570 sg13g2_dlygate4sd3_1
XFILLER_2_908 VPWR VGND sg13g2_decap_8
X_05167_ _01897_ _01894_ _01896_ _01612_ i_exotiny._0314_\[2\] VPWR VGND sg13g2_a22oi_1
XFILLER_104_825 VPWR VGND sg13g2_decap_8
Xhold787 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[30\]
+ VPWR VGND net2614 sg13g2_dlygate4sd3_1
Xhold776 _00293_ VPWR VGND net2603 sg13g2_dlygate4sd3_1
Xhold765 i_exotiny._0022_\[3\] VPWR VGND net2592 sg13g2_dlygate4sd3_1
XFILLER_103_346 VPWR VGND sg13g2_decap_8
X_09225__754 VPWR VGND net754 sg13g2_tiehi
Xhold798 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[17\]
+ VPWR VGND net2625 sg13g2_dlygate4sd3_1
X_05098_ _01825_ _01826_ _01827_ _01828_ VPWR VGND sg13g2_or3_1
XFILLER_39_37 VPWR VGND sg13g2_fill_2
Xhold1410 _01128_ VPWR VGND net3237 sg13g2_dlygate4sd3_1
X_08926_ net1476 VGND VPWR net2760 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[24\]
+ clknet_leaf_65_clk_regs sg13g2_dfrbpq_1
Xhold1443 i_exotiny._0026_\[2\] VPWR VGND net3270 sg13g2_dlygate4sd3_1
XFILLER_58_945 VPWR VGND sg13g2_fill_2
Xhold1421 _00738_ VPWR VGND net3248 sg13g2_dlygate4sd3_1
X_08857_ net1549 VGND VPWR net2712 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[24\]
+ clknet_leaf_185_clk_regs sg13g2_dfrbpq_1
Xhold1432 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[16\]
+ VPWR VGND net3259 sg13g2_dlygate4sd3_1
Xhold1454 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[6\]
+ VPWR VGND net3281 sg13g2_dlygate4sd3_1
Xhold1465 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[11\]
+ VPWR VGND net3292 sg13g2_dlygate4sd3_1
Xhold1476 _00310_ VPWR VGND net3303 sg13g2_dlygate4sd3_1
X_07808_ net2862 net2733 net892 _01287_ VPWR VGND sg13g2_mux2_1
X_08449__231 VPWR VGND net231 sg13g2_tiehi
XFILLER_45_606 VPWR VGND sg13g2_decap_4
Xhold1498 _00503_ VPWR VGND net3325 sg13g2_dlygate4sd3_1
Xhold1487 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[4\]
+ VPWR VGND net3314 sg13g2_dlygate4sd3_1
X_08788_ net1620 VGND VPWR net2118 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[19\]
+ clknet_leaf_164_clk_regs sg13g2_dfrbpq_1
XFILLER_44_127 VPWR VGND sg13g2_fill_1
X_07739_ net1227 _01576_ net1118 _03205_ VPWR VGND sg13g2_nor3_1
X_09156__826 VPWR VGND net826 sg13g2_tiehi
X_09232__747 VPWR VGND net747 sg13g2_tiehi
X_08456__224 VPWR VGND net224 sg13g2_tiehi
XFILLER_105_0 VPWR VGND sg13g2_fill_2
X_08645__1332 VPWR VGND net1752 sg13g2_tiehi
X_09163__819 VPWR VGND net819 sg13g2_tiehi
XFILLER_106_195 VPWR VGND sg13g2_decap_8
XFILLER_95_517 VPWR VGND sg13g2_fill_2
XFILLER_1_985 VPWR VGND sg13g2_decap_8
Xhold70 i_exotiny.i_wb_spi.dat_rx_r\[11\] VPWR VGND net1897 sg13g2_dlygate4sd3_1
Xhold81 _00029_ VPWR VGND net1908 sg13g2_dlygate4sd3_1
Xhold92 _00053_ VPWR VGND net1919 sg13g2_dlygate4sd3_1
XFILLER_36_628 VPWR VGND sg13g2_decap_8
XFILLER_75_274 VPWR VGND sg13g2_fill_1
X_08463__217 VPWR VGND net217 sg13g2_tiehi
XFILLER_90_277 VPWR VGND sg13g2_fill_1
XFILLER_44_661 VPWR VGND sg13g2_fill_2
X_08183__494 VPWR VGND net494 sg13g2_tiehi
XFILLER_12_591 VPWR VGND sg13g2_fill_2
X_06070_ _02517_ net1262 _02475_ VPWR VGND sg13g2_nand2_2
XFILLER_6_63 VPWR VGND sg13g2_fill_2
X_05021_ _01753_ net1238 net1240 VPWR VGND sg13g2_nand2_2
XFILLER_99_856 VPWR VGND sg13g2_decap_8
XFILLER_98_355 VPWR VGND sg13g2_decap_8
X_06972_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[14\]
+ net2329 net1020 _00745_ VPWR VGND sg13g2_mux2_1
X_05923_ net886 i_exotiny._0019_\[0\] _02478_ _02480_ VPWR VGND sg13g2_mux2_1
XFILLER_20_0 VPWR VGND sg13g2_fill_2
X_08711_ net1697 VGND VPWR _00769_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[6\]
+ clknet_leaf_116_clk_regs sg13g2_dfrbpq_1
Xfanout1090 net1091 net1090 VPWR VGND sg13g2_buf_8
X_08190__487 VPWR VGND net487 sg13g2_tiehi
X_08642_ net1755 VGND VPWR net2849 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[11\]
+ clknet_leaf_145_clk_regs sg13g2_dfrbpq_1
XFILLER_66_274 VPWR VGND sg13g2_fill_2
XFILLER_26_127 VPWR VGND sg13g2_fill_2
X_05854_ _02443_ i_exotiny._0352_ _01470_ VPWR VGND sg13g2_nand2_1
X_05785_ net3709 VPWR _00074_ VGND _02390_ _02406_ sg13g2_o21ai_1
X_04805_ _01551_ net1127 VPWR VGND net1233 sg13g2_nand2b_2
X_08573_ net58 VGND VPWR _00646_ i_exotiny._0314_\[18\] clknet_leaf_166_clk_regs sg13g2_dfrbpq_1
X_04736_ _01492_ net3724 _01491_ VPWR VGND sg13g2_nand2_1
X_07524_ _03106_ VPWR _03121_ VGND _01500_ _01872_ sg13g2_o21ai_1
XFILLER_50_631 VPWR VGND sg13g2_fill_2
X_07455_ VGND VPWR net3609 net1080 _03093_ _03077_ sg13g2_a21oi_1
X_04667_ net1250 net1252 net1253 _01428_ VPWR VGND sg13g2_nor3_2
X_06406_ net1071 net3759 _02589_ _00513_ VPWR VGND sg13g2_a21o_1
X_08723__1265 VPWR VGND net1685 sg13g2_tiehi
X_07386_ net2026 net1078 _03040_ VPWR VGND sg13g2_nor2_1
X_06337_ _02561_ net3147 net1033 _00472_ VPWR VGND sg13g2_mux2_1
X_09125_ net857 VGND VPWR net3139 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[13\]
+ clknet_leaf_154_clk_regs sg13g2_dfrbpq_1
X_09056_ net1346 VGND VPWR net1971 i_exotiny.i_rstctl.cnt\[6\] clknet_leaf_40_clk_regs
+ sg13g2_dfrbpq_1
X_06268_ net3179 i_exotiny._0016_\[0\] net942 _00411_ VPWR VGND sg13g2_mux2_1
X_08007_ net688 VGND VPWR _00088_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[8\]
+ clknet_leaf_62_clk_regs sg13g2_dfrbpq_1
X_05219_ _01947_ _01632_ i_exotiny._0022_\[1\] _01628_ i_exotiny._0037_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold540 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[21\]
+ VPWR VGND net2367 sg13g2_dlygate4sd3_1
X_06199_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[11\]
+ net3495 net947 _00354_ VPWR VGND sg13g2_mux2_1
Xhold551 _00186_ VPWR VGND net2378 sg13g2_dlygate4sd3_1
Xhold562 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[25\]
+ VPWR VGND net2389 sg13g2_dlygate4sd3_1
Xhold584 _00795_ VPWR VGND net2411 sg13g2_dlygate4sd3_1
Xhold573 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[29\]
+ VPWR VGND net2400 sg13g2_dlygate4sd3_1
Xhold595 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[18\]
+ VPWR VGND net2422 sg13g2_dlygate4sd3_1
XFILLER_106_31 VPWR VGND sg13g2_decap_8
XFILLER_104_699 VPWR VGND sg13g2_decap_8
XFILLER_103_143 VPWR VGND sg13g2_decap_8
X_08945__1037 VPWR VGND net1457 sg13g2_tiehi
X_08909_ net1493 VGND VPWR net2468 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[7\]
+ clknet_leaf_113_clk_regs sg13g2_dfrbpq_1
XFILLER_106_97 VPWR VGND sg13g2_decap_8
XFILLER_100_861 VPWR VGND sg13g2_decap_8
XFILLER_85_561 VPWR VGND sg13g2_fill_2
XFILLER_57_230 VPWR VGND sg13g2_fill_1
Xhold1240 _01359_ VPWR VGND net3067 sg13g2_dlygate4sd3_1
Xhold1251 _00793_ VPWR VGND net3078 sg13g2_dlygate4sd3_1
XFILLER_72_211 VPWR VGND sg13g2_fill_1
Xhold1262 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[13\]
+ VPWR VGND net3089 sg13g2_dlygate4sd3_1
Xhold1273 _00739_ VPWR VGND net3100 sg13g2_dlygate4sd3_1
Xhold1284 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[4\]
+ VPWR VGND net3111 sg13g2_dlygate4sd3_1
Xhold1295 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[18\]
+ VPWR VGND net3122 sg13g2_dlygate4sd3_1
XFILLER_40_163 VPWR VGND sg13g2_fill_2
XFILLER_41_697 VPWR VGND sg13g2_decap_4
X_09030__952 VPWR VGND net1372 sg13g2_tiehi
X_09261__239 VPWR VGND net239 sg13g2_tiehi
XFILLER_95_314 VPWR VGND sg13g2_decap_8
X_09208__771 VPWR VGND net771 sg13g2_tiehi
XFILLER_1_782 VPWR VGND sg13g2_decap_8
XFILLER_95_369 VPWR VGND sg13g2_decap_8
X_08801__1187 VPWR VGND net1607 sg13g2_tiehi
X_09139__843 VPWR VGND net843 sg13g2_tiehi
X_05570_ _02250_ i_exotiny._0315_\[8\] _02249_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_141 VPWR VGND sg13g2_fill_2
X_07240_ net2467 net3049 net1005 _00963_ VPWR VGND sg13g2_mux2_1
X_09215__764 VPWR VGND net764 sg13g2_tiehi
X_07171_ i_exotiny._0036_\[0\] net886 _02947_ _02949_ VPWR VGND sg13g2_mux2_1
X_06122_ net2979 net2539 net1046 _00291_ VPWR VGND sg13g2_mux2_1
XFILLER_106_909 VPWR VGND sg13g2_decap_8
X_09146__836 VPWR VGND net836 sg13g2_tiehi
X_06053_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[25\]
+ net2391 net961 _00238_ VPWR VGND sg13g2_mux2_1
X_05004_ _01734_ _01735_ _01736_ VPWR VGND sg13g2_and2_1
XFILLER_99_697 VPWR VGND sg13g2_fill_2
X_09222__757 VPWR VGND net757 sg13g2_tiehi
XFILLER_95_870 VPWR VGND sg13g2_decap_8
XFILLER_74_509 VPWR VGND sg13g2_fill_1
X_06955_ net2575 _02921_ net927 _00730_ VPWR VGND sg13g2_mux2_1
XFILLER_39_241 VPWR VGND sg13g2_fill_1
X_05906_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[11\]
+ net2903 net973 _00123_ VPWR VGND sg13g2_mux2_1
X_06886_ VGND VPWR net1094 _02891_ _00690_ _02892_ sg13g2_a21oi_1
X_08625_ net1770 VGND VPWR _00697_ i_exotiny.i_rstctl.wdg_res_n clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_2
X_07943__87 VPWR VGND net87 sg13g2_tiehi
X_05837_ _02426_ _01497_ net1224 _01431_ _01427_ VPWR VGND sg13g2_a22oi_1
X_08446__234 VPWR VGND net234 sg13g2_tiehi
X_08556_ net100 VGND VPWR net3604 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[1\].i_hadd.a_i
+ clknet_leaf_5_clk_regs sg13g2_dfrbpq_2
X_05768_ _02396_ i_exotiny._2034_\[3\] net1127 VPWR VGND sg13g2_nand2_1
X_09153__829 VPWR VGND net829 sg13g2_tiehi
X_07507_ net2841 i_exotiny._0315_\[20\] net901 _01090_ VPWR VGND sg13g2_mux2_1
X_05699_ net1982 net1059 _02345_ VPWR VGND sg13g2_nor2_1
X_08487_ net193 VGND VPWR _00561_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[7\]
+ clknet_leaf_110_clk_regs sg13g2_dfrbpq_1
X_04719_ _01477_ net3819 _01475_ VPWR VGND sg13g2_nand2_1
X_07438_ _03081_ _03008_ net1149 net1209 net3535 VPWR VGND sg13g2_a22oi_1
XFILLER_11_859 VPWR VGND sg13g2_fill_2
X_07369_ VGND VPWR net1077 _03027_ _01038_ _03024_ sg13g2_a21oi_1
X_09108_ net1294 VGND VPWR net3086 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[28\]
+ clknet_leaf_141_clk_regs sg13g2_dfrbpq_1
X_09039_ net1363 VGND VPWR _01097_ i_exotiny._0315_\[27\] clknet_leaf_181_clk_regs
+ sg13g2_dfrbpq_1
X_08453__227 VPWR VGND net227 sg13g2_tiehi
Xhold370 _00497_ VPWR VGND net2197 sg13g2_dlygate4sd3_1
Xhold381 _00178_ VPWR VGND net2208 sg13g2_dlygate4sd3_1
XFILLER_105_986 VPWR VGND sg13g2_decap_8
XFILLER_104_474 VPWR VGND sg13g2_decap_8
Xhold392 _00323_ VPWR VGND net2219 sg13g2_dlygate4sd3_1
XFILLER_81_1015 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_179_clk_regs clknet_5_1__leaf_clk_regs clknet_leaf_179_clk_regs VPWR
+ VGND sg13g2_buf_8
Xclkbuf_leaf_108_clk_regs clknet_5_28__leaf_clk_regs clknet_leaf_108_clk_regs VPWR
+ VGND sg13g2_buf_8
Xfanout883 net884 net883 VPWR VGND sg13g2_buf_8
Xfanout894 net895 net894 VPWR VGND sg13g2_buf_8
Xfanout872 _02472_ net872 VPWR VGND sg13g2_buf_8
X_07991__132 VPWR VGND net132 sg13g2_tiehi
Xhold1081 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[20\]
+ VPWR VGND net2908 sg13g2_dlygate4sd3_1
Xhold1070 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[29\]
+ VPWR VGND net2897 sg13g2_dlygate4sd3_1
Xhold1092 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[24\]
+ VPWR VGND net2919 sg13g2_dlygate4sd3_1
XFILLER_34_907 VPWR VGND sg13g2_fill_1
XFILLER_73_564 VPWR VGND sg13g2_fill_2
XFILLER_60_236 VPWR VGND sg13g2_fill_1
X_08145__540 VPWR VGND net540 sg13g2_tiehi
X_08819__1169 VPWR VGND net1589 sg13g2_tiehi
X_08180__497 VPWR VGND net497 sg13g2_tiehi
XFILLER_6_885 VPWR VGND sg13g2_decap_4
XFILLER_5_395 VPWR VGND sg13g2_fill_2
XFILLER_69_826 VPWR VGND sg13g2_fill_2
XFILLER_96_656 VPWR VGND sg13g2_fill_1
XFILLER_95_111 VPWR VGND sg13g2_fill_1
X_06740_ VGND VPWR _02767_ _02769_ _02770_ net1130 sg13g2_a21oi_1
XFILLER_3_1026 VPWR VGND sg13g2_fill_2
X_08545__111 VPWR VGND net111 sg13g2_tiehi
X_06671_ _02691_ VPWR _02709_ VGND _02688_ _02708_ sg13g2_o21ai_1
X_08410_ net275 VGND VPWR _00484_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[9\]
+ clknet_leaf_89_clk_regs sg13g2_dfrbpq_1
X_05622_ VGND VPWR net1061 _02287_ _00031_ _02285_ sg13g2_a21oi_1
XFILLER_91_383 VPWR VGND sg13g2_fill_1
X_08341_ net337 VGND VPWR net2386 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[11\]
+ clknet_leaf_98_clk_regs sg13g2_dfrbpq_1
X_07948__708 VPWR VGND net708 sg13g2_tiehi
X_05553_ VGND VPWR _01523_ _02236_ _02237_ _01553_ sg13g2_a21oi_1
X_08272_ net406 VGND VPWR _00353_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[6\]
+ clknet_leaf_100_clk_regs sg13g2_dfrbpq_1
X_05484_ _02183_ net1283 _01512_ VPWR VGND sg13g2_nand2_1
Xclkbuf_5_18__f_clk_regs clknet_4_9_0_clk_regs clknet_5_18__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07223_ i_exotiny.i_wb_spi.dat_rx_r\[19\] net3644 net1086 _00948_ VPWR VGND sg13g2_mux2_1
XFILLER_106_706 VPWR VGND sg13g2_decap_8
X_07154_ net3107 net2858 net1009 _00902_ VPWR VGND sg13g2_mux2_1
X_06105_ net2400 _02522_ net955 _00279_ VPWR VGND sg13g2_mux2_1
X_08552__104 VPWR VGND net104 sg13g2_tiehi
X_07085_ net2144 net3197 net913 _00840_ VPWR VGND sg13g2_mux2_1
XFILLER_105_249 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_6_clk_regs clknet_5_2__leaf_clk_regs clknet_leaf_6_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06036_ net2464 net2637 net964 _00221_ VPWR VGND sg13g2_mux2_1
XFILLER_102_923 VPWR VGND sg13g2_decap_8
XFILLER_99_472 VPWR VGND sg13g2_decap_8
XFILLER_101_422 VPWR VGND sg13g2_decap_8
X_08559__92 VPWR VGND net92 sg13g2_tiehi
X_07975__116 VPWR VGND net116 sg13g2_tiehi
X_07987_ net128 VGND VPWR net2062 i_exotiny._0369_\[11\] clknet_leaf_165_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_101_499 VPWR VGND sg13g2_decap_8
XFILLER_86_177 VPWR VGND sg13g2_fill_1
X_06938_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[18\]
+ net2278 net925 _00717_ VPWR VGND sg13g2_mux2_1
X_06869_ i_exotiny._0369_\[28\] net1189 _02878_ VPWR VGND sg13g2_nor2_1
X_09020__962 VPWR VGND net1382 sg13g2_tiehi
X_08608_ net1788 VGND VPWR net3718 i_exotiny._1617_\[0\] clknet_leaf_23_clk_regs sg13g2_dfrbpq_2
X_08895__1087 VPWR VGND net1507 sg13g2_tiehi
X_08539_ net141 VGND VPWR _00613_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[27\]
+ clknet_leaf_182_clk_regs sg13g2_dfrbpq_1
XFILLER_3_844 VPWR VGND sg13g2_decap_8
X_09129__853 VPWR VGND net853 sg13g2_tiehi
XFILLER_105_783 VPWR VGND sg13g2_decap_8
XFILLER_104_271 VPWR VGND sg13g2_decap_8
X_08682__1306 VPWR VGND net1726 sg13g2_tiehi
XFILLER_34_737 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_76_clk_regs clknet_5_26__leaf_clk_regs clknet_leaf_76_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_61_578 VPWR VGND sg13g2_fill_1
X_09136__846 VPWR VGND net846 sg13g2_tiehi
XFILLER_61_589 VPWR VGND sg13g2_fill_1
X_09212__767 VPWR VGND net767 sg13g2_tiehi
X_08940__1042 VPWR VGND net1462 sg13g2_tiehi
XFILLER_97_954 VPWR VGND sg13g2_decap_8
X_07910_ net738 VGND VPWR net1904 i_exotiny._1924_\[3\] clknet_leaf_31_clk_regs sg13g2_dfrbpq_1
X_08890_ net1512 VGND VPWR net3645 i_exotiny.i_wb_spi.dat_rx_r\[20\] clknet_leaf_63_clk_regs
+ sg13g2_dfrbpq_1
X_09143__839 VPWR VGND net839 sg13g2_tiehi
Xhold1817 i_exotiny.i_wb_spi.dat_rx_r\[20\] VPWR VGND net3644 sg13g2_dlygate4sd3_1
XFILLER_25_1027 VPWR VGND sg13g2_fill_2
X_07841_ net2347 net3254 net986 _01314_ VPWR VGND sg13g2_mux2_1
Xhold1806 _00660_ VPWR VGND net3633 sg13g2_dlygate4sd3_1
X_07772_ net3007 net3290 net990 _01257_ VPWR VGND sg13g2_mux2_1
Xhold1839 i_exotiny.i_wdg_top.o_wb_dat\[2\] VPWR VGND net3666 sg13g2_dlygate4sd3_1
Xhold1828 i_exotiny.i_wb_spi.dat_rx_r\[19\] VPWR VGND net3655 sg13g2_dlygate4sd3_1
X_06723_ _02756_ _02719_ net3808 net1068 net3567 VPWR VGND sg13g2_a22oi_1
XFILLER_56_339 VPWR VGND sg13g2_fill_1
X_04984_ net1242 net1250 _01716_ VPWR VGND sg13g2_nor2_1
XFILLER_83_158 VPWR VGND sg13g2_fill_1
X_06654_ _02694_ VPWR _02695_ VGND _02690_ _02692_ sg13g2_o21ai_1
X_05605_ _01397_ _01366_ net1116 _02275_ VPWR VGND sg13g2_mux2_1
X_06585_ net1199 _02645_ _02646_ _00635_ VPWR VGND sg13g2_nor3_1
X_08324_ net354 VGND VPWR _00405_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[26\]
+ clknet_leaf_73_clk_regs sg13g2_dfrbpq_1
X_05536_ _02223_ net3706 VPWR VGND net1272 sg13g2_nand2b_2
X_08255_ net422 VGND VPWR _00336_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[22\]
+ clknet_leaf_49_clk_regs sg13g2_dfrbpq_1
X_05467_ VPWR VGND i_exotiny._1616_\[3\] _02172_ _02146_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s2wto.u_bit_field.i_sw_write_data[0]
+ _02173_ _02145_ sg13g2_a221oi_1
X_05398_ _01401_ _02110_ _02114_ VPWR VGND sg13g2_and2_1
X_07206_ net1933 net2105 net1089 _00938_ VPWR VGND sg13g2_mux2_1
X_08186_ net491 VGND VPWR net3280 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[17\]
+ clknet_leaf_111_clk_regs sg13g2_dfrbpq_1
XFILLER_106_503 VPWR VGND sg13g2_decap_8
X_07137_ net1286 net1866 _00887_ VPWR VGND sg13g2_and2_1
X_08760__1228 VPWR VGND net1648 sg13g2_tiehi
XFILLER_4_619 VPWR VGND sg13g2_fill_1
X_07068_ net3065 net874 _02934_ _02939_ VPWR VGND sg13g2_mux2_1
XFILLER_102_731 VPWR VGND sg13g2_decap_8
X_06019_ _00019_ net1103 _02504_ VPWR VGND sg13g2_nor2_1
XFILLER_87_420 VPWR VGND sg13g2_fill_1
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_88_965 VPWR VGND sg13g2_decap_8
XFILLER_102_797 VPWR VGND sg13g2_decap_8
XFILLER_101_296 VPWR VGND sg13g2_decap_8
XFILLER_28_531 VPWR VGND sg13g2_decap_8
XFILLER_90_607 VPWR VGND sg13g2_fill_1
XFILLER_15_225 VPWR VGND sg13g2_fill_1
XFILLER_43_523 VPWR VGND sg13g2_fill_2
XFILLER_90_89 VPWR VGND sg13g2_fill_2
XFILLER_8_958 VPWR VGND sg13g2_decap_8
X_08142__543 VPWR VGND net543 sg13g2_tiehi
XFILLER_7_479 VPWR VGND sg13g2_fill_2
X_08736__1252 VPWR VGND net1672 sg13g2_tiehi
XFILLER_97_206 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_123_clk_regs clknet_5_22__leaf_clk_regs clknet_leaf_123_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_94_913 VPWR VGND sg13g2_decap_8
XFILLER_78_442 VPWR VGND sg13g2_fill_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_94_1025 VPWR VGND sg13g2_decap_4
X_08958__1024 VPWR VGND net1444 sg13g2_tiehi
X_06370_ net2576 net3053 net1028 _00500_ VPWR VGND sg13g2_mux2_1
XFILLER_9_96 VPWR VGND sg13g2_fill_1
XFILLER_9_74 VPWR VGND sg13g2_fill_2
X_05321_ VPWR VGND net1110 _02042_ _02014_ i_exotiny._0550_ _02045_ _01829_ sg13g2_a221oi_1
X_08040_ net654 VGND VPWR net2553 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[9\]
+ clknet_leaf_55_clk_regs sg13g2_dfrbpq_1
X_05252_ _01976_ _01977_ _01972_ _01978_ VPWR VGND sg13g2_nand3_1
Xhold903 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[25\]
+ VPWR VGND net2730 sg13g2_dlygate4sd3_1
Xhold914 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[28\]
+ VPWR VGND net2741 sg13g2_dlygate4sd3_1
XFILLER_50_0 VPWR VGND sg13g2_decap_8
Xhold936 _00290_ VPWR VGND net2763 sg13g2_dlygate4sd3_1
Xhold925 _01279_ VPWR VGND net2752 sg13g2_dlygate4sd3_1
X_05183_ _01908_ _01910_ _01911_ VPWR VGND sg13g2_and2_1
Xhold947 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[26\]
+ VPWR VGND net2774 sg13g2_dlygate4sd3_1
Xhold958 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[16\]
+ VPWR VGND net2785 sg13g2_dlygate4sd3_1
Xhold969 _00246_ VPWR VGND net2796 sg13g2_dlygate4sd3_1
X_09010__972 VPWR VGND net1392 sg13g2_tiehi
XFILLER_103_528 VPWR VGND sg13g2_decap_8
X_08942_ net1460 VGND VPWR _01000_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[8\]
+ clknet_leaf_75_clk_regs sg13g2_dfrbpq_1
Xhold1614 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[18\]
+ VPWR VGND net3441 sg13g2_dlygate4sd3_1
Xhold1603 i_exotiny._2025_\[6\] VPWR VGND net3430 sg13g2_dlygate4sd3_1
X_08873_ net1529 VGND VPWR net3575 i_exotiny.i_wb_spi.dat_rx_r\[3\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_1
Xhold1625 i_exotiny._0032_\[3\] VPWR VGND net3452 sg13g2_dlygate4sd3_1
XFILLER_96_294 VPWR VGND sg13g2_decap_8
Xhold1669 _00354_ VPWR VGND net3496 sg13g2_dlygate4sd3_1
XFILLER_56_125 VPWR VGND sg13g2_fill_2
Xhold1647 _01341_ VPWR VGND net3474 sg13g2_dlygate4sd3_1
Xhold1658 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[5\]
+ VPWR VGND net3485 sg13g2_dlygate4sd3_1
Xhold1636 _00638_ VPWR VGND net3463 sg13g2_dlygate4sd3_1
X_07824_ net2134 i_exotiny._0022_\[0\] net987 _01297_ VPWR VGND sg13g2_mux2_1
X_07755_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[11\]
+ net2460 net990 _01240_ VPWR VGND sg13g2_mux2_1
XFILLER_72_607 VPWR VGND sg13g2_fill_1
X_04967_ _01363_ _01692_ _01699_ VPWR VGND sg13g2_nor2_1
X_06706_ VGND VPWR _02739_ _02740_ _02741_ _02721_ sg13g2_a21oi_1
X_07686_ net2194 net2978 net998 _01188_ VPWR VGND sg13g2_mux2_1
X_04898_ net1256 _01617_ _01623_ _01630_ VPWR VGND sg13g2_nor3_2
X_06637_ net2008 net1159 _02681_ VPWR VGND sg13g2_nor2_1
X_08814__1174 VPWR VGND net1594 sg13g2_tiehi
X_09119__863 VPWR VGND net863 sg13g2_tiehi
X_06568_ i_exotiny._0314_\[2\] net1162 _02635_ VPWR VGND sg13g2_nor2_1
X_08307_ net371 VGND VPWR _00388_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[9\]
+ clknet_leaf_83_clk_regs sg13g2_dfrbpq_1
X_06499_ net2341 net2659 net1026 _00580_ VPWR VGND sg13g2_mux2_1
X_09287_ net1825 VGND VPWR net2212 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[13\]
+ clknet_leaf_179_clk_regs sg13g2_dfrbpq_1
X_05519_ _02209_ net2997 net1069 VPWR VGND sg13g2_nand2_1
X_08238_ net439 VGND VPWR net3278 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[5\]
+ clknet_leaf_57_clk_regs sg13g2_dfrbpq_1
XFILLER_20_261 VPWR VGND sg13g2_fill_1
XFILLER_106_300 VPWR VGND sg13g2_decap_8
XFILLER_5_917 VPWR VGND sg13g2_decap_8
X_08169_ net508 VGND VPWR _00250_ i_exotiny._0038_\[0\] clknet_leaf_110_clk_regs sg13g2_dfrbpq_2
X_09272__77 VPWR VGND net77 sg13g2_tiehi
XFILLER_106_377 VPWR VGND sg13g2_decap_8
X_09126__856 VPWR VGND net856 sg13g2_tiehi
XFILLER_47_103 VPWR VGND sg13g2_fill_2
XFILLER_87_283 VPWR VGND sg13g2_fill_2
XFILLER_91_938 VPWR VGND sg13g2_decap_8
XFILLER_18_72 VPWR VGND sg13g2_fill_1
XFILLER_18_83 VPWR VGND sg13g2_fill_2
X_09172__810 VPWR VGND net810 sg13g2_tiehi
XFILLER_44_865 VPWR VGND sg13g2_fill_2
XFILLER_70_172 VPWR VGND sg13g2_fill_2
X_09133__849 VPWR VGND net849 sg13g2_tiehi
XFILLER_102_1007 VPWR VGND sg13g2_decap_8
XFILLER_12_784 VPWR VGND sg13g2_fill_1
XFILLER_79_751 VPWR VGND sg13g2_fill_2
XFILLER_3_493 VPWR VGND sg13g2_fill_1
Xfanout1250 net1251 net1250 VPWR VGND sg13g2_buf_8
X_08890__1092 VPWR VGND net1512 sg13g2_tiehi
Xfanout1283 net1285 net1283 VPWR VGND sg13g2_buf_8
Xfanout1261 net3804 net1261 VPWR VGND sg13g2_buf_8
Xfanout1272 net1274 net1272 VPWR VGND sg13g2_buf_8
X_05870_ _02456_ VPWR _02457_ VGND _01911_ _02267_ sg13g2_o21ai_1
X_04821_ net1867 net1868 net1865 net1839 _01561_ VPWR VGND sg13g2_nor4_1
Xclkbuf_leaf_91_clk_regs clknet_5_31__leaf_clk_regs clknet_leaf_91_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_93_275 VPWR VGND sg13g2_decap_8
X_04752_ _01502_ _01505_ _01501_ _00001_ VPWR VGND sg13g2_nand3_1
X_07540_ VGND VPWR _03128_ _03132_ _01104_ net1196 sg13g2_a21oi_1
Xclkbuf_leaf_20_clk_regs clknet_5_12__leaf_clk_regs clknet_leaf_20_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_90_982 VPWR VGND sg13g2_decap_8
X_07471_ _03103_ VPWR _01064_ VGND _02988_ _03094_ sg13g2_o21ai_1
X_04683_ net3832 net3824 net3834 _01443_ VPWR VGND sg13g2_nand3_1
X_06422_ _02600_ _02601_ _00517_ VPWR VGND sg13g2_nor2_1
XFILLER_22_537 VPWR VGND sg13g2_fill_2
X_09210_ net769 VGND VPWR net3228 i_exotiny._0023_\[0\] clknet_leaf_129_clk_regs sg13g2_dfrbpq_2
X_06353_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[12\]
+ net2929 net1029 _00483_ VPWR VGND sg13g2_mux2_1
X_09141_ net841 VGND VPWR _01196_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[29\]
+ clknet_leaf_154_clk_regs sg13g2_dfrbpq_1
X_09072_ net1330 VGND VPWR net1892 i_exotiny.i_wdg_top.clk_div_inst.cnt\[12\] clknet_5_11__leaf_clk_regs
+ sg13g2_dfrbpq_1
X_05304_ _02030_ _01631_ i_exotiny._0027_\[0\] _01624_ i_exotiny._0040_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_06284_ net2698 net2507 net942 _00427_ VPWR VGND sg13g2_mux2_1
X_08023_ net671 VGND VPWR _00104_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[24\]
+ clknet_leaf_63_clk_regs sg13g2_dfrbpq_1
Xhold711 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[9\]
+ VPWR VGND net2538 sg13g2_dlygate4sd3_1
Xhold700 _01187_ VPWR VGND net2527 sg13g2_dlygate4sd3_1
X_05235_ _01963_ _01654_ i_exotiny._0020_\[1\] _01634_ i_exotiny._0013_\[1\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_104_804 VPWR VGND sg13g2_decap_8
Xhold722 _00803_ VPWR VGND net2549 sg13g2_dlygate4sd3_1
Xhold755 _01247_ VPWR VGND net2582 sg13g2_dlygate4sd3_1
Xhold733 _01260_ VPWR VGND net2560 sg13g2_dlygate4sd3_1
Xhold744 _02914_ VPWR VGND net2571 sg13g2_dlygate4sd3_1
X_05166_ _01612_ _01895_ _01896_ VPWR VGND sg13g2_nor2_1
XFILLER_103_325 VPWR VGND sg13g2_decap_8
Xhold766 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[25\]
+ VPWR VGND net2593 sg13g2_dlygate4sd3_1
Xhold788 _00990_ VPWR VGND net2615 sg13g2_dlygate4sd3_1
Xhold777 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[13\]
+ VPWR VGND net2604 sg13g2_dlygate4sd3_1
Xhold799 _01282_ VPWR VGND net2626 sg13g2_dlygate4sd3_1
X_05097_ _01826_ _01827_ net37 VPWR VGND sg13g2_nor2_1
X_08925_ net1477 VGND VPWR _00983_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[23\]
+ clknet_leaf_66_clk_regs sg13g2_dfrbpq_1
Xhold1400 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[4\]
+ VPWR VGND net3227 sg13g2_dlygate4sd3_1
Xhold1433 i_exotiny._0014_\[0\] VPWR VGND net3260 sg13g2_dlygate4sd3_1
X_08856_ net1550 VGND VPWR net2443 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[23\]
+ clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
Xhold1422 i_exotiny._0023_\[3\] VPWR VGND net3249 sg13g2_dlygate4sd3_1
Xhold1411 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[20\]
+ VPWR VGND net3238 sg13g2_dlygate4sd3_1
Xhold1477 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[28\]
+ VPWR VGND net3304 sg13g2_dlygate4sd3_1
XFILLER_85_787 VPWR VGND sg13g2_fill_1
Xhold1455 i_exotiny._0018_\[2\] VPWR VGND net3282 sg13g2_dlygate4sd3_1
Xhold1444 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[14\]
+ VPWR VGND net3271 sg13g2_dlygate4sd3_1
Xhold1466 _01272_ VPWR VGND net3293 sg13g2_dlygate4sd3_1
X_07807_ net2850 net2680 net894 _01286_ VPWR VGND sg13g2_mux2_1
Xhold1499 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.genblk7.g_value.r_value[0]
+ VPWR VGND net3326 sg13g2_dlygate4sd3_1
Xhold1488 _00964_ VPWR VGND net3315 sg13g2_dlygate4sd3_1
X_08787_ net1621 VGND VPWR _00845_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[18\]
+ clknet_leaf_169_clk_regs sg13g2_dfrbpq_1
XFILLER_38_670 VPWR VGND sg13g2_fill_2
XFILLER_38_692 VPWR VGND sg13g2_fill_1
XFILLER_44_106 VPWR VGND sg13g2_decap_8
X_05999_ net2669 net2898 net1048 _00201_ VPWR VGND sg13g2_mux2_1
XFILLER_53_640 VPWR VGND sg13g2_decap_8
X_07738_ _03204_ net2547 net996 _01230_ VPWR VGND sg13g2_mux2_1
XFILLER_52_161 VPWR VGND sg13g2_fill_2
X_07669_ net2182 net2980 net1000 _01171_ VPWR VGND sg13g2_mux2_1
X_10680_ gpo net33 VPWR VGND sg13g2_buf_1
XFILLER_52_183 VPWR VGND sg13g2_fill_2
XFILLER_13_537 VPWR VGND sg13g2_fill_2
XFILLER_84_1024 VPWR VGND sg13g2_decap_4
XFILLER_5_769 VPWR VGND sg13g2_decap_8
XFILLER_106_174 VPWR VGND sg13g2_decap_8
XFILLER_103_881 VPWR VGND sg13g2_decap_8
XFILLER_1_964 VPWR VGND sg13g2_decap_8
XFILLER_76_743 VPWR VGND sg13g2_fill_1
Xhold60 _01118_ VPWR VGND net1887 sg13g2_dlygate4sd3_1
Xhold82 i_exotiny._1924_\[11\] VPWR VGND net1909 sg13g2_dlygate4sd3_1
Xhold71 _00940_ VPWR VGND net1898 sg13g2_dlygate4sd3_1
XFILLER_63_404 VPWR VGND sg13g2_fill_1
Xhold93 i_exotiny._1924_\[25\] VPWR VGND net1920 sg13g2_dlygate4sd3_1
XFILLER_29_681 VPWR VGND sg13g2_fill_1
XFILLER_90_234 VPWR VGND sg13g2_fill_1
XFILLER_28_191 VPWR VGND sg13g2_fill_1
XFILLER_16_364 VPWR VGND sg13g2_fill_2
X_09000__982 VPWR VGND net1402 sg13g2_tiehi
X_05020_ _01751_ VPWR _01752_ VGND _01745_ _01749_ sg13g2_o21ai_1
XFILLER_99_835 VPWR VGND sg13g2_decap_8
XFILLER_98_334 VPWR VGND sg13g2_decap_8
XFILLER_101_829 VPWR VGND sg13g2_decap_8
X_06971_ net2988 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[17\]
+ net1018 _00744_ VPWR VGND sg13g2_mux2_1
X_09109__873 VPWR VGND net1293 sg13g2_tiehi
XFILLER_100_339 VPWR VGND sg13g2_decap_8
X_05922_ net2668 net2430 net973 _00139_ VPWR VGND sg13g2_mux2_1
X_08710_ net1698 VGND VPWR net2090 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[5\]
+ clknet_leaf_121_clk_regs sg13g2_dfrbpq_1
XFILLER_67_754 VPWR VGND sg13g2_fill_1
Xfanout1091 net1092 net1091 VPWR VGND sg13g2_buf_8
XFILLER_66_253 VPWR VGND sg13g2_fill_1
X_08641_ net1756 VGND VPWR net2784 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[10\]
+ clknet_leaf_149_clk_regs sg13g2_dfrbpq_1
XFILLER_13_0 VPWR VGND sg13g2_fill_1
X_05853_ _02442_ _02440_ _02441_ VPWR VGND sg13g2_nand2_1
Xfanout1080 net1084 net1080 VPWR VGND sg13g2_buf_8
X_04804_ i_exotiny._0315_\[2\] _01549_ _01550_ VPWR VGND sg13g2_nor2_1
XFILLER_82_724 VPWR VGND sg13g2_fill_1
XFILLER_27_629 VPWR VGND sg13g2_fill_1
X_05784_ _02407_ net1126 _01373_ net1145 net3708 VPWR VGND sg13g2_a22oi_1
X_08572_ net60 VGND VPWR _00645_ i_exotiny._0314_\[17\] clknet_leaf_181_clk_regs sg13g2_dfrbpq_1
X_04735_ VGND VPWR _01488_ _01490_ _01491_ net1226 sg13g2_a21oi_1
XFILLER_23_813 VPWR VGND sg13g2_fill_1
X_07523_ net3470 _02462_ _03120_ VPWR VGND sg13g2_nor2_1
X_07454_ _03092_ net1148 _03028_ net1207 net3415 VPWR VGND sg13g2_a22oi_1
X_04666_ net1252 net1253 _01427_ VPWR VGND sg13g2_nor2_2
XFILLER_50_654 VPWR VGND sg13g2_decap_8
X_06405_ _02219_ _02587_ _02588_ _02589_ VPWR VGND sg13g2_nor3_1
XFILLER_50_698 VPWR VGND sg13g2_decap_4
X_07385_ VGND VPWR net1077 _03038_ _01042_ _03039_ sg13g2_a21oi_1
X_09116__866 VPWR VGND net866 sg13g2_tiehi
X_06336_ i_exotiny._0014_\[1\] net882 _02558_ _02561_ VPWR VGND sg13g2_mux2_1
X_09124_ net858 VGND VPWR net2421 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[12\]
+ clknet_leaf_152_clk_regs sg13g2_dfrbpq_1
X_09055_ net1347 VGND VPWR _01110_ i_exotiny.i_rstctl.cnt\[5\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_2
X_08299__379 VPWR VGND net379 sg13g2_tiehi
X_06267_ VGND VPWR net1140 _02552_ _02553_ net1166 sg13g2_a21oi_1
X_08555__102 VPWR VGND net102 sg13g2_tiehi
Xhold530 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[20\]
+ VPWR VGND net2357 sg13g2_dlygate4sd3_1
X_08006_ net689 VGND VPWR _00087_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[7\]
+ clknet_leaf_62_clk_regs sg13g2_dfrbpq_1
X_05218_ _01946_ _01637_ i_exotiny._0024_\[1\] _01636_ i_exotiny._0019_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold541 _00432_ VPWR VGND net2368 sg13g2_dlygate4sd3_1
X_06198_ net2427 net2565 net948 _00353_ VPWR VGND sg13g2_mux2_1
Xhold563 _00307_ VPWR VGND net2390 sg13g2_dlygate4sd3_1
Xhold552 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[29\]
+ VPWR VGND net2379 sg13g2_dlygate4sd3_1
XFILLER_103_122 VPWR VGND sg13g2_decap_8
Xhold574 _00275_ VPWR VGND net2401 sg13g2_dlygate4sd3_1
Xhold585 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[24\]
+ VPWR VGND net2412 sg13g2_dlygate4sd3_1
X_09162__820 VPWR VGND net820 sg13g2_tiehi
Xhold596 _01213_ VPWR VGND net2423 sg13g2_dlygate4sd3_1
X_05149_ VPWR VGND i_exotiny._0039_\[2\] _01878_ _01651_ i_exotiny._0034_\[2\] _01879_
+ _01619_ sg13g2_a221oi_1
XFILLER_104_678 VPWR VGND sg13g2_decap_4
XFILLER_106_76 VPWR VGND sg13g2_decap_8
XFILLER_103_199 VPWR VGND sg13g2_decap_8
X_08908_ net1494 VGND VPWR net2362 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[6\]
+ clknet_leaf_65_clk_regs sg13g2_dfrbpq_1
X_09123__859 VPWR VGND net859 sg13g2_tiehi
XFILLER_100_840 VPWR VGND sg13g2_decap_8
Xhold1230 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[10\]
+ VPWR VGND net3057 sg13g2_dlygate4sd3_1
Xhold1241 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[20\]
+ VPWR VGND net3068 sg13g2_dlygate4sd3_1
Xhold1252 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[17\]
+ VPWR VGND net3079 sg13g2_dlygate4sd3_1
Xhold1274 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[21\]
+ VPWR VGND net3101 sg13g2_dlygate4sd3_1
X_08839_ net1567 VGND VPWR _00897_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[6\]
+ clknet_leaf_185_clk_regs sg13g2_dfrbpq_1
Xhold1263 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[20\]
+ VPWR VGND net3090 sg13g2_dlygate4sd3_1
Xhold1285 _00282_ VPWR VGND net3112 sg13g2_dlygate4sd3_1
Xhold1296 i_exotiny._0031_\[0\] VPWR VGND net3123 sg13g2_dlygate4sd3_1
XFILLER_40_153 VPWR VGND sg13g2_fill_1
XFILLER_5_544 VPWR VGND sg13g2_decap_4
X_09302__1113 VPWR VGND net1533 sg13g2_tiehi
XFILLER_1_761 VPWR VGND sg13g2_decap_8
XFILLER_0_260 VPWR VGND sg13g2_fill_2
X_08773__1215 VPWR VGND net1635 sg13g2_tiehi
X_08599__1377 VPWR VGND net1797 sg13g2_tiehi
XFILLER_37_949 VPWR VGND sg13g2_fill_1
XFILLER_45_993 VPWR VGND sg13g2_fill_2
Xclkbuf_5_17__f_clk_regs clknet_4_8_0_clk_regs clknet_5_17__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
X_07170_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[31\]
+ net2956 net1008 _00918_ VPWR VGND sg13g2_mux2_1
X_06121_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[12\]
+ net2762 net1043 _00290_ VPWR VGND sg13g2_mux2_1
X_06052_ net2257 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[20\]
+ net964 _00237_ VPWR VGND sg13g2_mux2_1
XFILLER_99_610 VPWR VGND sg13g2_fill_1
X_05003_ _01735_ _01366_ _01712_ VPWR VGND sg13g2_nand2_1
XFILLER_98_197 VPWR VGND sg13g2_fill_1
X_06954_ net2720 net873 _02916_ _02921_ VPWR VGND sg13g2_mux2_1
X_05905_ net2817 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[14\]
+ net973 _00122_ VPWR VGND sg13g2_mux2_1
X_06885_ net3672 net1094 _02892_ VPWR VGND sg13g2_nor2_1
X_08624_ net1772 VGND VPWR net3467 i_exotiny._1586_ clknet_leaf_38_clk_regs sg13g2_dfrbpq_2
X_05836_ VGND VPWR net1242 _01458_ _02425_ _01817_ sg13g2_a21oi_1
X_05767_ _02395_ VPWR _00068_ VGND net1143 _02394_ sg13g2_o21ai_1
XFILLER_54_267 VPWR VGND sg13g2_fill_1
X_08555_ net102 VGND VPWR net3494 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_pc.genblk3\[0\].i_hadd.a_i
+ clknet_leaf_4_clk_regs sg13g2_dfrbpq_2
XFILLER_63_790 VPWR VGND sg13g2_fill_2
X_07506_ net3185 net3625 net904 _01089_ VPWR VGND sg13g2_mux2_1
X_08486_ net194 VGND VPWR net2531 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[6\]
+ clknet_leaf_93_clk_regs sg13g2_dfrbpq_1
X_05698_ VGND VPWR net1061 _02344_ _00050_ _02342_ sg13g2_a21oi_1
X_04718_ VPWR _01476_ _01475_ VGND sg13g2_inv_1
X_04649_ VPWR _01411_ i_exotiny.i_wb_spi.dat_rx_r\[8\] VGND sg13g2_inv_1
X_07437_ _03080_ VPWR _01053_ VGND net1082 _03079_ sg13g2_o21ai_1
X_07368_ _03027_ _03025_ _03026_ net1212 net1996 VPWR VGND sg13g2_a22oi_1
X_09107_ net1295 VGND VPWR _01162_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[27\]
+ clknet_leaf_144_clk_regs sg13g2_dfrbpq_1
X_06319_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[17\]
+ net2650 net1034 _00456_ VPWR VGND sg13g2_mux2_1
X_07299_ net2662 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[28\]
+ net909 _01016_ VPWR VGND sg13g2_mux2_1
X_09038_ net1364 VGND VPWR _01096_ i_exotiny._0315_\[26\] clknet_leaf_179_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_105_965 VPWR VGND sg13g2_decap_8
Xhold371 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[17\]
+ VPWR VGND net2198 sg13g2_dlygate4sd3_1
Xhold360 _01136_ VPWR VGND net2187 sg13g2_dlygate4sd3_1
XFILLER_104_453 VPWR VGND sg13g2_decap_8
Xhold382 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[31\]
+ VPWR VGND net2209 sg13g2_dlygate4sd3_1
Xhold393 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[16\]
+ VPWR VGND net2220 sg13g2_dlygate4sd3_1
Xfanout884 net885 net884 VPWR VGND sg13g2_buf_8
Xfanout873 net875 net873 VPWR VGND sg13g2_buf_8
XFILLER_85_370 VPWR VGND sg13g2_fill_1
Xhold1060 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[27\]
+ VPWR VGND net2887 sg13g2_dlygate4sd3_1
XFILLER_19_938 VPWR VGND sg13g2_fill_1
Xfanout895 _03217_ net895 VPWR VGND sg13g2_buf_8
Xhold1093 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[10\]
+ VPWR VGND net2920 sg13g2_dlygate4sd3_1
X_08169__508 VPWR VGND net508 sg13g2_tiehi
Xhold1082 _00751_ VPWR VGND net2909 sg13g2_dlygate4sd3_1
Xhold1071 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[29\]
+ VPWR VGND net2898 sg13g2_dlygate4sd3_1
XFILLER_45_245 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_148_clk_regs clknet_5_16__leaf_clk_regs clknet_leaf_148_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08827__1161 VPWR VGND net1581 sg13g2_tiehi
XFILLER_6_864 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
X_09106__876 VPWR VGND net1296 sg13g2_tiehi
XFILLER_3_1005 VPWR VGND sg13g2_decap_8
X_06670_ _02263_ net3390 _02708_ VPWR VGND sg13g2_xor2_1
X_05621_ VGND VPWR i_exotiny._1612_\[1\] net1120 _02287_ _02286_ sg13g2_a21oi_1
X_08289__389 VPWR VGND net389 sg13g2_tiehi
XFILLER_51_215 VPWR VGND sg13g2_fill_2
X_08340_ net338 VGND VPWR net2776 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[10\]
+ clknet_leaf_95_clk_regs sg13g2_dfrbpq_1
X_05552_ i_exotiny._0315_\[21\] i_exotiny._0314_\[21\] net1272 _02236_ VPWR VGND sg13g2_mux2_1
X_08271_ net407 VGND VPWR _00352_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[5\]
+ clknet_leaf_106_clk_regs sg13g2_dfrbpq_1
X_09152__830 VPWR VGND net830 sg13g2_tiehi
X_05483_ net1076 VPWR i_exotiny._1611_\[7\] VGND _02175_ _02182_ sg13g2_o21ai_1
X_07222_ net1937 net3655 net1087 _00947_ VPWR VGND sg13g2_mux2_1
X_07153_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[14\]
+ net2787 net1010 _00901_ VPWR VGND sg13g2_mux2_1
X_09113__869 VPWR VGND net869 sg13g2_tiehi
X_06104_ net2791 net883 _02519_ _02522_ VPWR VGND sg13g2_mux2_1
X_07084_ net3076 net2967 net913 _00839_ VPWR VGND sg13g2_mux2_1
XFILLER_105_228 VPWR VGND sg13g2_decap_8
X_06035_ net2513 i_exotiny._0025_\[3\] net963 _00220_ VPWR VGND sg13g2_mux2_1
XFILLER_102_902 VPWR VGND sg13g2_decap_8
XFILLER_99_451 VPWR VGND sg13g2_decap_8
XFILLER_101_401 VPWR VGND sg13g2_decap_8
XFILLER_102_979 VPWR VGND sg13g2_decap_8
X_07986_ net127 VGND VPWR net3308 i_exotiny._0369_\[10\] clknet_leaf_166_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_101_478 VPWR VGND sg13g2_decap_8
X_06937_ net2265 net2503 net924 _00716_ VPWR VGND sg13g2_mux2_1
XFILLER_27_201 VPWR VGND sg13g2_fill_1
XFILLER_82_340 VPWR VGND sg13g2_fill_1
X_08607_ net1789 VGND VPWR _00679_ i_exotiny._1614_\[3\] clknet_leaf_23_clk_regs sg13g2_dfrbpq_2
X_06868_ VGND VPWR net1095 _02876_ _00687_ _02877_ sg13g2_a21oi_1
XFILLER_82_373 VPWR VGND sg13g2_fill_2
X_05819_ net2597 net2540 net1054 _00091_ VPWR VGND sg13g2_mux2_1
X_06799_ VGND VPWR net3717 net1130 _02820_ net3734 sg13g2_a21oi_1
X_08538_ net142 VGND VPWR net2966 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[26\]
+ clknet_leaf_184_clk_regs sg13g2_dfrbpq_1
X_08469_ net211 VGND VPWR _00543_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[21\]
+ clknet_leaf_163_clk_regs sg13g2_dfrbpq_1
XFILLER_12_74 VPWR VGND sg13g2_fill_2
XFILLER_3_823 VPWR VGND sg13g2_decap_8
XFILLER_105_762 VPWR VGND sg13g2_decap_8
XFILLER_104_250 VPWR VGND sg13g2_decap_8
Xhold190 _00465_ VPWR VGND net2017 sg13g2_dlygate4sd3_1
XFILLER_78_657 VPWR VGND sg13g2_fill_2
X_08565__74 VPWR VGND net74 sg13g2_tiehi
XFILLER_101_990 VPWR VGND sg13g2_decap_8
X_08628__743 VPWR VGND net743 sg13g2_tiehi
XFILLER_37_82 VPWR VGND sg13g2_fill_2
XFILLER_37_93 VPWR VGND sg13g2_fill_1
XFILLER_73_373 VPWR VGND sg13g2_fill_2
XFILLER_33_204 VPWR VGND sg13g2_fill_1
XFILLER_18_1002 VPWR VGND sg13g2_fill_1
XFILLER_30_966 VPWR VGND sg13g2_fill_2
XFILLER_30_999 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_45_clk_regs clknet_5_11__leaf_clk_regs clknet_leaf_45_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_97_933 VPWR VGND sg13g2_decap_8
Xhold1807 i_exotiny.i_wb_spi.state_r\[0\] VPWR VGND net3634 sg13g2_dlygate4sd3_1
Xhold1818 _00948_ VPWR VGND net3645 sg13g2_dlygate4sd3_1
X_07840_ net2469 net3259 net986 _01313_ VPWR VGND sg13g2_mux2_1
X_07771_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[27\]
+ net2519 net990 _01256_ VPWR VGND sg13g2_mux2_1
Xhold1829 i_exotiny.i_wb_regs.spi_auto_cs_o VPWR VGND net3656 sg13g2_dlygate4sd3_1
XFILLER_65_852 VPWR VGND sg13g2_fill_1
X_06722_ VPWR VGND net7 _02754_ _02747_ net3785 _02755_ net1182 sg13g2_a221oi_1
XFILLER_49_392 VPWR VGND sg13g2_fill_2
XFILLER_49_381 VPWR VGND sg13g2_fill_2
X_04983_ VGND VPWR _01361_ _01712_ _01715_ _01714_ sg13g2_a21oi_1
XFILLER_65_885 VPWR VGND sg13g2_fill_1
XFILLER_64_362 VPWR VGND sg13g2_fill_2
XFILLER_64_351 VPWR VGND sg13g2_fill_1
X_08850__1136 VPWR VGND net1556 sg13g2_tiehi
XFILLER_37_576 VPWR VGND sg13g2_decap_4
XFILLER_52_513 VPWR VGND sg13g2_fill_1
X_06653_ i_exotiny._0352_ net1153 _02693_ _02694_ VPWR VGND sg13g2_nor3_1
X_05604_ net1978 net1060 _02274_ VPWR VGND sg13g2_nor2_1
X_06584_ net3517 net1155 _02646_ VPWR VGND sg13g2_nor2_1
X_08323_ net355 VGND VPWR _00404_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[25\]
+ clknet_leaf_72_clk_regs sg13g2_dfrbpq_1
X_05535_ _02222_ net2864 net1272 VPWR VGND sg13g2_nand2_1
X_09269__83 VPWR VGND net83 sg13g2_tiehi
X_08254_ net423 VGND VPWR net2227 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[21\]
+ clknet_leaf_57_clk_regs sg13g2_dfrbpq_1
X_05466_ _02170_ _02171_ _02169_ _02172_ VPWR VGND sg13g2_nand3_1
X_09284__53 VPWR VGND net53 sg13g2_tiehi
X_05397_ _01401_ _02110_ _02113_ VPWR VGND sg13g2_nor2_1
X_07205_ _02964_ VPWR _00937_ VGND _01411_ net1088 sg13g2_o21ai_1
X_08185_ net492 VGND VPWR _00266_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[16\]
+ clknet_leaf_110_clk_regs sg13g2_dfrbpq_1
X_07136_ net1286 net1838 _00886_ VPWR VGND sg13g2_and2_1
X_07067_ _02938_ net2313 net1017 _00825_ VPWR VGND sg13g2_mux2_1
X_08594__1382 VPWR VGND net1802 sg13g2_tiehi
XFILLER_106_559 VPWR VGND sg13g2_decap_8
X_06018_ VGND VPWR net2042 net1103 _00211_ _02503_ sg13g2_a21oi_1
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_102_776 VPWR VGND sg13g2_decap_8
XFILLER_101_275 VPWR VGND sg13g2_decap_8
XFILLER_59_178 VPWR VGND sg13g2_fill_2
X_07969_ net1175 VGND VPWR net1889 i_exotiny.i_wdg_top.o_wb_dat\[10\] clknet_leaf_33_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_56_830 VPWR VGND sg13g2_fill_2
XFILLER_23_270 VPWR VGND sg13g2_fill_2
XFILLER_8_937 VPWR VGND sg13g2_decap_8
XFILLER_12_988 VPWR VGND sg13g2_decap_8
X_08279__399 VPWR VGND net399 sg13g2_tiehi
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_105_592 VPWR VGND sg13g2_decap_8
XFILLER_66_616 VPWR VGND sg13g2_fill_1
X_08631__1346 VPWR VGND net1766 sg13g2_tiehi
Xclkbuf_leaf_163_clk_regs clknet_5_5__leaf_clk_regs clknet_leaf_163_clk_regs VPWR
+ VGND sg13g2_buf_8
X_09142__840 VPWR VGND net840 sg13g2_tiehi
XFILLER_94_969 VPWR VGND sg13g2_decap_8
XFILLER_62_800 VPWR VGND sg13g2_fill_2
X_09103__879 VPWR VGND net1299 sg13g2_tiehi
XFILLER_0_1008 VPWR VGND sg13g2_decap_8
XFILLER_94_1004 VPWR VGND sg13g2_decap_8
XFILLER_74_671 VPWR VGND sg13g2_fill_2
XFILLER_62_833 VPWR VGND sg13g2_fill_2
XFILLER_22_708 VPWR VGND sg13g2_fill_2
XFILLER_34_546 VPWR VGND sg13g2_fill_2
XFILLER_14_292 VPWR VGND sg13g2_fill_2
X_05320_ _02043_ _02044_ net38 VPWR VGND sg13g2_nor2_2
XFILLER_30_774 VPWR VGND sg13g2_fill_1
X_05251_ _01831_ _01974_ _01975_ _01977_ VPWR VGND sg13g2_or3_1
X_09266__97 VPWR VGND net97 sg13g2_tiehi
Xhold904 _00468_ VPWR VGND net2731 sg13g2_dlygate4sd3_1
X_05182_ _01905_ _01907_ _01910_ VPWR VGND _01900_ sg13g2_nand3b_1
Xhold937 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[22\]
+ VPWR VGND net2764 sg13g2_dlygate4sd3_1
Xhold915 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[29\]
+ VPWR VGND net2742 sg13g2_dlygate4sd3_1
Xhold926 i_exotiny._0043_\[1\] VPWR VGND net2753 sg13g2_dlygate4sd3_1
XFILLER_103_507 VPWR VGND sg13g2_decap_8
Xhold948 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[14\]
+ VPWR VGND net2775 sg13g2_dlygate4sd3_1
Xhold959 _01151_ VPWR VGND net2786 sg13g2_dlygate4sd3_1
X_08941_ net1461 VGND VPWR _00999_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[7\]
+ clknet_leaf_51_clk_regs sg13g2_dfrbpq_1
X_08872_ net1530 VGND VPWR net3577 i_exotiny.i_wb_spi.dat_rx_r\[2\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_96_273 VPWR VGND sg13g2_decap_8
Xhold1604 i_exotiny._1902_\[6\] VPWR VGND net3431 sg13g2_dlygate4sd3_1
Xhold1626 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[23\].i_reg.reg_r\[26\]
+ VPWR VGND net3453 sg13g2_dlygate4sd3_1
Xhold1615 i_exotiny._0037_\[3\] VPWR VGND net3442 sg13g2_dlygate4sd3_1
X_07823_ VGND VPWR net1138 _03222_ _03223_ net1168 sg13g2_a21oi_1
Xhold1637 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[26\]
+ VPWR VGND net3464 sg13g2_dlygate4sd3_1
Xhold1648 i_exotiny._0314_\[10\] VPWR VGND net3475 sg13g2_dlygate4sd3_1
Xhold1659 _00218_ VPWR VGND net3486 sg13g2_dlygate4sd3_1
X_07754_ net3057 net3256 net988 _01239_ VPWR VGND sg13g2_mux2_1
XFILLER_56_148 VPWR VGND sg13g2_fill_2
X_04966_ _01698_ i_exotiny.i_fazyrv_top.i_fazyrv_core.cntrl_icyc\[2\] _01696_ VPWR
+ VGND sg13g2_nand2_1
XFILLER_93_991 VPWR VGND sg13g2_decap_8
XFILLER_53_811 VPWR VGND sg13g2_fill_2
X_06705_ _02740_ _02723_ net17 _02593_ i_exotiny._2025_\[5\] VPWR VGND sg13g2_a22oi_1
X_07685_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[20\]
+ net2526 net1000 _01187_ VPWR VGND sg13g2_mux2_1
X_06636_ net1195 _02679_ _02680_ _00652_ VPWR VGND sg13g2_nor3_1
X_08786__1202 VPWR VGND net1622 sg13g2_tiehi
X_04897_ _01629_ i_exotiny._0037_\[3\] _01628_ VPWR VGND sg13g2_nand2_1
X_06567_ net1200 _02633_ _02634_ _00629_ VPWR VGND sg13g2_nor3_1
X_08306_ net372 VGND VPWR net2987 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[8\]
+ clknet_leaf_82_clk_regs sg13g2_dfrbpq_1
X_06498_ net2532 net2583 net1025 _00579_ VPWR VGND sg13g2_mux2_1
X_09286_ net42 VGND VPWR net3474 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[12\]
+ clknet_leaf_175_clk_regs sg13g2_dfrbpq_1
X_05518_ _02206_ VPWR i_exotiny._1611_\[19\] VGND net1075 _02208_ sg13g2_o21ai_1
X_08237_ net440 VGND VPWR _00318_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[4\]
+ clknet_leaf_55_clk_regs sg13g2_dfrbpq_1
X_05449_ _02157_ _02146_ i_exotiny._1616_\[1\] _02145_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_rvd1.u_bit_field.i_sw_write_data[0]
+ VPWR VGND sg13g2_a22oi_1
X_08168_ net510 VGND VPWR net2141 i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_spm_d.repl_r
+ clknet_leaf_8_clk_regs sg13g2_dfrbpq_1
XFILLER_106_356 VPWR VGND sg13g2_decap_8
X_07119_ net1288 net1853 _00869_ VPWR VGND sg13g2_and2_1
X_08099_ net595 VGND VPWR _00180_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[4\]
+ clknet_leaf_124_clk_regs sg13g2_dfrbpq_1
XFILLER_83_490 VPWR VGND sg13g2_fill_1
XFILLER_31_549 VPWR VGND sg13g2_fill_2
XFILLER_15_1016 VPWR VGND sg13g2_decap_8
XFILLER_15_1027 VPWR VGND sg13g2_fill_2
X_08649__1328 VPWR VGND net1748 sg13g2_tiehi
XFILLER_98_516 VPWR VGND sg13g2_decap_8
XFILLER_4_995 VPWR VGND sg13g2_decap_8
Xfanout1240 net1241 net1240 VPWR VGND sg13g2_buf_8
Xfanout1262 net3144 net1262 VPWR VGND sg13g2_buf_8
Xfanout1273 net1274 net1273 VPWR VGND sg13g2_buf_8
Xfanout1251 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[4\]
+ net1251 VPWR VGND sg13g2_buf_2
X_04820_ net1852 net1845 net1856 net1843 _01560_ VPWR VGND sg13g2_nor4_1
Xfanout1284 net1285 net1284 VPWR VGND sg13g2_buf_1
XFILLER_81_416 VPWR VGND sg13g2_fill_1
XFILLER_75_991 VPWR VGND sg13g2_fill_1
X_08907__1075 VPWR VGND net1495 sg13g2_tiehi
X_04751_ VPWR VGND net1273 net1196 net1212 net1201 _01505_ _01454_ sg13g2_a221oi_1
XFILLER_90_961 VPWR VGND sg13g2_decap_8
XFILLER_34_376 VPWR VGND sg13g2_fill_2
X_07470_ _03076_ VPWR _03103_ VGND _02997_ net1147 sg13g2_o21ai_1
X_04682_ _01442_ net3832 net3824 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_60_clk_regs clknet_5_13__leaf_clk_regs clknet_leaf_60_clk_regs VPWR VGND
+ sg13g2_buf_8
X_06421_ net1282 VPWR _02601_ VGND net3561 net3689 sg13g2_o21ai_1
X_06352_ net2269 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[7\]
+ net1030 _00482_ VPWR VGND sg13g2_mux2_1
X_09140_ net842 VGND VPWR net2977 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[28\]
+ clknet_leaf_158_clk_regs sg13g2_dfrbpq_1
X_09071_ net1331 VGND VPWR _01126_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[11\] clknet_leaf_46_clk_regs
+ sg13g2_dfrbpq_1
X_06283_ net3405 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[15\]
+ net943 _00426_ VPWR VGND sg13g2_mux2_1
X_05303_ _02029_ _01649_ i_exotiny._0042_\[0\] _01625_ i_exotiny._0030_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_08022_ net672 VGND VPWR _00103_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[23\]
+ clknet_leaf_60_clk_regs sg13g2_dfrbpq_1
Xhold701 i_exotiny._1924_\[24\] VPWR VGND net2528 sg13g2_dlygate4sd3_1
Xhold712 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[9\]
+ VPWR VGND net2539 sg13g2_dlygate4sd3_1
X_05234_ _01962_ _01655_ i_exotiny._0026_\[1\] _01646_ i_exotiny._0017_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold745 _00698_ VPWR VGND net2572 sg13g2_dlygate4sd3_1
Xhold734 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[28\]
+ VPWR VGND net2561 sg13g2_dlygate4sd3_1
Xhold723 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[10\]
+ VPWR VGND net2550 sg13g2_dlygate4sd3_1
X_05165_ i_exotiny._0036_\[2\] _01644_ _01895_ VPWR VGND sg13g2_nor2_1
XFILLER_103_304 VPWR VGND sg13g2_decap_8
Xhold756 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[25\]
+ VPWR VGND net2583 sg13g2_dlygate4sd3_1
Xhold767 _00271_ VPWR VGND net2594 sg13g2_dlygate4sd3_1
Xhold778 _00226_ VPWR VGND net2605 sg13g2_dlygate4sd3_1
X_05096_ _01607_ _01676_ _01827_ VPWR VGND sg13g2_and2_1
Xhold789 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[22\]
+ VPWR VGND net2616 sg13g2_dlygate4sd3_1
X_08924_ net1478 VGND VPWR _00982_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[22\]
+ clknet_leaf_64_clk_regs sg13g2_dfrbpq_1
Xhold1401 _01265_ VPWR VGND net3228 sg13g2_dlygate4sd3_1
Xhold1434 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[5\]
+ VPWR VGND net3261 sg13g2_dlygate4sd3_1
XFILLER_69_295 VPWR VGND sg13g2_fill_1
Xhold1423 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[18\]
+ VPWR VGND net3250 sg13g2_dlygate4sd3_1
X_08855_ net1551 VGND VPWR _00913_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[22\]
+ clknet_leaf_186_clk_regs sg13g2_dfrbpq_1
Xhold1412 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[30\]
+ VPWR VGND net3239 sg13g2_dlygate4sd3_1
Xhold1456 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[20\]
+ VPWR VGND net3283 sg13g2_dlygate4sd3_1
Xhold1467 i_exotiny._0027_\[0\] VPWR VGND net3294 sg13g2_dlygate4sd3_1
Xhold1445 _01209_ VPWR VGND net3272 sg13g2_dlygate4sd3_1
X_08786_ net1622 VGND VPWR net2159 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[17\]
+ clknet_leaf_168_clk_regs sg13g2_dfrbpq_1
X_07806_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[20\]
+ net3225 net895 _01285_ VPWR VGND sg13g2_mux2_1
Xhold1478 _00823_ VPWR VGND net3305 sg13g2_dlygate4sd3_1
Xhold1489 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[17\]
+ VPWR VGND net3316 sg13g2_dlygate4sd3_1
X_05998_ net2754 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[28\]
+ net1050 _00200_ VPWR VGND sg13g2_mux2_1
X_07737_ net3459 net872 _03199_ _03204_ VPWR VGND sg13g2_mux2_1
X_04949_ VGND VPWR net1242 net1184 _01681_ _01466_ sg13g2_a21oi_1
X_07668_ i_exotiny._0030_\[3\] net2633 net1001 _01170_ VPWR VGND sg13g2_mux2_1
X_07599_ net1205 net1878 _03170_ _01125_ VPWR VGND sg13g2_nor3_1
X_06619_ i_exotiny._0314_\[19\] net1160 _02669_ VPWR VGND sg13g2_nor2_1
X_09132__850 VPWR VGND net850 sg13g2_tiehi
X_09269_ net83 VGND VPWR net2268 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[27\]
+ clknet_leaf_130_clk_regs sg13g2_dfrbpq_1
XFILLER_105_2 VPWR VGND sg13g2_fill_1
XFILLER_84_1003 VPWR VGND sg13g2_decap_8
XFILLER_106_153 VPWR VGND sg13g2_decap_8
XFILLER_96_34 VPWR VGND sg13g2_fill_1
XFILLER_1_943 VPWR VGND sg13g2_decap_8
XFILLER_103_860 VPWR VGND sg13g2_decap_8
Xhold50 i_exotiny.i_wdg_top.clk_div_inst.cnt\[10\] VPWR VGND net1877 sg13g2_dlygate4sd3_1
XFILLER_29_61 VPWR VGND sg13g2_fill_2
XFILLER_102_392 VPWR VGND sg13g2_decap_8
Xhold61 _00020_ VPWR VGND net1888 sg13g2_dlygate4sd3_1
Xhold83 _00036_ VPWR VGND net1910 sg13g2_dlygate4sd3_1
Xhold72 i_exotiny._1924_\[29\] VPWR VGND net1899 sg13g2_dlygate4sd3_1
Xhold94 _00050_ VPWR VGND net1921 sg13g2_dlygate4sd3_1
Xhold1990 i_exotiny._1618_\[2\] VPWR VGND net3817 sg13g2_dlygate4sd3_1
XFILLER_35_118 VPWR VGND sg13g2_fill_1
XFILLER_43_140 VPWR VGND sg13g2_fill_2
XFILLER_44_663 VPWR VGND sg13g2_fill_1
Xclkbuf_5_16__f_clk_regs clknet_4_8_0_clk_regs clknet_5_16__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_12_593 VPWR VGND sg13g2_fill_1
XFILLER_8_542 VPWR VGND sg13g2_fill_2
XFILLER_98_313 VPWR VGND sg13g2_decap_8
XFILLER_4_792 VPWR VGND sg13g2_decap_8
XFILLER_101_808 VPWR VGND sg13g2_decap_8
X_06970_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[12\]
+ net2722 net1021 _00743_ VPWR VGND sg13g2_mux2_1
XFILLER_100_318 VPWR VGND sg13g2_decap_8
X_05921_ net2481 net2509 net974 _00138_ VPWR VGND sg13g2_mux2_1
XFILLER_6_1025 VPWR VGND sg13g2_decap_4
XFILLER_20_2 VPWR VGND sg13g2_fill_1
Xfanout1092 net1093 net1092 VPWR VGND sg13g2_buf_8
Xfanout1070 _02181_ net1070 VPWR VGND sg13g2_buf_8
X_08640_ net1757 VGND VPWR net2857 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[9\]
+ clknet_leaf_147_clk_regs sg13g2_dfrbpq_1
X_05852_ _02055_ _02069_ _02439_ _02441_ VPWR VGND sg13g2_or3_1
Xfanout1081 net1084 net1081 VPWR VGND sg13g2_buf_2
X_04803_ _00026_ net1144 VPWR VGND sg13g2_inv_2
XFILLER_66_276 VPWR VGND sg13g2_fill_1
X_05783_ _02406_ i_exotiny._2034_\[8\] net1127 VPWR VGND sg13g2_nand2_1
X_08571_ net62 VGND VPWR net3359 i_exotiny._0314_\[16\] clknet_leaf_3_clk_regs sg13g2_dfrbpq_1
XFILLER_19_181 VPWR VGND sg13g2_fill_1
XFILLER_26_129 VPWR VGND sg13g2_fill_1
X_04734_ net1231 net3713 _01383_ _01490_ VPWR VGND net1218 sg13g2_nand4_1
X_07522_ _03119_ net3377 net902 VPWR VGND sg13g2_nand2_1
X_07453_ _03091_ VPWR _01058_ VGND net1082 _03090_ sg13g2_o21ai_1
X_04665_ net3692 net3822 net3670 _01426_ VPWR VGND sg13g2_nor3_1
X_06404_ _01522_ _02586_ _02588_ VPWR VGND sg13g2_nor2_1
X_09123_ net859 VGND VPWR _01178_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[11\]
+ clknet_leaf_155_clk_regs sg13g2_dfrbpq_1
X_07384_ net1996 net1077 _03039_ VPWR VGND sg13g2_nor2_1
X_06335_ _02560_ net3223 net1034 _00471_ VPWR VGND sg13g2_mux2_1
X_09054_ net1348 VGND VPWR _01109_ i_exotiny.i_rstctl.cnt\[4\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_1
X_06266_ _02420_ _02509_ _02552_ VPWR VGND sg13g2_nor2_2
X_08005_ net690 VGND VPWR _00086_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[6\]
+ clknet_leaf_68_clk_regs sg13g2_dfrbpq_1
Xhold520 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[21\]
+ VPWR VGND net2347 sg13g2_dlygate4sd3_1
X_05217_ _01945_ _01920_ _01944_ net1108 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[1\]
+ VPWR VGND sg13g2_a22oi_1
Xhold531 _00128_ VPWR VGND net2358 sg13g2_dlygate4sd3_1
X_06197_ net2947 net2230 net945 _00352_ VPWR VGND sg13g2_mux2_1
Xhold542 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[21\]
+ VPWR VGND net2369 sg13g2_dlygate4sd3_1
Xhold553 _01224_ VPWR VGND net2380 sg13g2_dlygate4sd3_1
XFILLER_2_729 VPWR VGND sg13g2_fill_1
XFILLER_104_657 VPWR VGND sg13g2_decap_8
Xhold586 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[22\]
+ VPWR VGND net2413 sg13g2_dlygate4sd3_1
Xhold597 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[29\]
+ VPWR VGND net2424 sg13g2_dlygate4sd3_1
Xhold575 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[8\]
+ VPWR VGND net2402 sg13g2_dlygate4sd3_1
Xhold564 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[21\]
+ VPWR VGND net2391 sg13g2_dlygate4sd3_1
X_05148_ _01876_ _01877_ _01874_ _01878_ VPWR VGND sg13g2_nand3_1
X_05079_ VPWR VGND i_exotiny._0013_\[3\] _01810_ _01777_ i_exotiny._0014_\[3\] _01811_
+ _01760_ sg13g2_a221oi_1
XFILLER_106_55 VPWR VGND sg13g2_decap_8
XFILLER_103_178 VPWR VGND sg13g2_decap_8
XFILLER_58_722 VPWR VGND sg13g2_fill_1
X_08907_ net1495 VGND VPWR _00965_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[5\]
+ clknet_leaf_112_clk_regs sg13g2_dfrbpq_1
Xhold1231 _01243_ VPWR VGND net3058 sg13g2_dlygate4sd3_1
Xhold1220 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[31\]
+ VPWR VGND net3047 sg13g2_dlygate4sd3_1
XFILLER_85_563 VPWR VGND sg13g2_fill_1
XFILLER_85_530 VPWR VGND sg13g2_decap_4
Xhold1242 _00542_ VPWR VGND net3069 sg13g2_dlygate4sd3_1
X_08838_ net1568 VGND VPWR _00896_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[5\]
+ clknet_leaf_185_clk_regs sg13g2_dfrbpq_1
XFILLER_18_608 VPWR VGND sg13g2_fill_1
XFILLER_100_896 VPWR VGND sg13g2_decap_8
XFILLER_85_596 VPWR VGND sg13g2_fill_1
Xhold1275 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[7\]
+ VPWR VGND net3102 sg13g2_dlygate4sd3_1
XFILLER_58_788 VPWR VGND sg13g2_fill_2
XFILLER_57_265 VPWR VGND sg13g2_fill_1
Xhold1264 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[5\]
+ VPWR VGND net3091 sg13g2_dlygate4sd3_1
XFILLER_18_619 VPWR VGND sg13g2_fill_2
Xhold1253 i_exotiny._0015_\[2\] VPWR VGND net3080 sg13g2_dlygate4sd3_1
Xhold1286 i_exotiny._0315_\[26\] VPWR VGND net3113 sg13g2_dlygate4sd3_1
XFILLER_17_129 VPWR VGND sg13g2_fill_2
Xhold1297 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[9\]
+ VPWR VGND net3124 sg13g2_dlygate4sd3_1
X_08769_ net1639 VGND VPWR _00827_ i_exotiny._0015_\[0\] clknet_leaf_169_clk_regs
+ sg13g2_dfrbpq_2
XFILLER_26_674 VPWR VGND sg13g2_fill_1
X_08863__1123 VPWR VGND net1543 sg13g2_tiehi
XFILLER_40_165 VPWR VGND sg13g2_fill_1
XFILLER_31_40 VPWR VGND sg13g2_decap_8
Xoutput40 net40 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_1_740 VPWR VGND sg13g2_decap_8
XFILLER_95_349 VPWR VGND sg13g2_decap_8
XFILLER_31_143 VPWR VGND sg13g2_fill_1
XFILLER_82_4 VPWR VGND sg13g2_fill_1
XFILLER_72_91 VPWR VGND sg13g2_fill_1
XFILLER_9_862 VPWR VGND sg13g2_fill_2
XFILLER_8_361 VPWR VGND sg13g2_fill_2
X_06120_ net2632 net2115 net1046 _00289_ VPWR VGND sg13g2_mux2_1
X_06051_ net2018 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[19\]
+ net964 _00236_ VPWR VGND sg13g2_mux2_1
X_08298__380 VPWR VGND net380 sg13g2_tiehi
X_05002_ _01711_ VPWR _01734_ VGND _01732_ _01733_ sg13g2_o21ai_1
X_07957__700 VPWR VGND net700 sg13g2_tiehi
X_06953_ net2927 _02920_ net925 _00729_ VPWR VGND sg13g2_mux2_1
X_05904_ net2552 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[13\]
+ net972 _00121_ VPWR VGND sg13g2_mux2_1
X_06884_ VGND VPWR i_exotiny._1618_\[2\] net1128 _02891_ _02890_ sg13g2_a21oi_1
X_09122__860 VPWR VGND net860 sg13g2_tiehi
X_05835_ net2091 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[27\]
+ net1054 _00107_ VPWR VGND sg13g2_mux2_1
X_08623_ net1773 VGND VPWR _00695_ i_exotiny._1618_\[3\] clknet_leaf_8_clk_regs sg13g2_dfrbpq_2
X_05766_ _02395_ net1126 net2087 net1144 net3666 VPWR VGND sg13g2_a22oi_1
X_08554_ net103 VGND VPWR i_exotiny._1207_ i_exotiny.i_fazyrv_top.i_fazyrv_core.i_fazyrv_alu.cmp_r
+ clknet_leaf_2_clk_regs sg13g2_dfrbpq_1
X_08644__1333 VPWR VGND net1753 sg13g2_tiehi
X_07505_ i_exotiny._0315_\[22\] net3549 net905 _01088_ VPWR VGND sg13g2_mux2_1
X_04717_ _01443_ _01474_ _01475_ VPWR VGND sg13g2_nor2_1
X_08485_ net195 VGND VPWR net2984 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[7\].i_reg.reg_r\[5\]
+ clknet_leaf_70_clk_regs sg13g2_dfrbpq_1
X_05697_ VGND VPWR i_exotiny._1619_\[0\] net1117 _02344_ _02343_ sg13g2_a21oi_1
X_04648_ VPWR _01410_ net1968 VGND sg13g2_inv_1
XFILLER_10_316 VPWR VGND sg13g2_fill_2
X_07436_ VGND VPWR net3541 net1082 _03080_ _03077_ sg13g2_a21oi_1
X_07367_ i_exotiny._0369_\[25\] net1213 _03026_ VPWR VGND sg13g2_and2_1
X_06318_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[11\].i_reg.reg_r\[16\]
+ net2325 net1035 _00455_ VPWR VGND sg13g2_mux2_1
X_09106_ net1296 VGND VPWR _01161_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[26\]
+ clknet_leaf_143_clk_regs sg13g2_dfrbpq_1
X_07298_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[23\]
+ net3471 net911 _01015_ VPWR VGND sg13g2_mux2_1
X_09037_ net1365 VGND VPWR net3221 i_exotiny._0315_\[25\] clknet_leaf_1_clk_regs sg13g2_dfrbpq_1
X_06249_ net3357 net2939 net1038 _00398_ VPWR VGND sg13g2_mux2_1
XFILLER_105_944 VPWR VGND sg13g2_decap_8
XFILLER_104_432 VPWR VGND sg13g2_decap_8
Xhold361 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[15\]
+ VPWR VGND net2188 sg13g2_dlygate4sd3_1
Xhold350 _01186_ VPWR VGND net2177 sg13g2_dlygate4sd3_1
X_08902__1080 VPWR VGND net1500 sg13g2_tiehi
Xhold372 _00904_ VPWR VGND net2199 sg13g2_dlygate4sd3_1
Xhold383 _01194_ VPWR VGND net2210 sg13g2_dlygate4sd3_1
Xhold394 _00233_ VPWR VGND net2221 sg13g2_dlygate4sd3_1
X_09260__241 VPWR VGND net241 sg13g2_tiehi
Xfanout874 net875 net874 VPWR VGND sg13g2_buf_8
Xfanout885 _02454_ net885 VPWR VGND sg13g2_buf_8
Xhold1050 _00567_ VPWR VGND net2877 sg13g2_dlygate4sd3_1
Xfanout896 net897 net896 VPWR VGND sg13g2_buf_8
Xhold1094 _00801_ VPWR VGND net2921 sg13g2_dlygate4sd3_1
Xhold1061 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[29\]
+ VPWR VGND net2888 sg13g2_dlygate4sd3_1
Xhold1083 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[29\]
+ VPWR VGND net2910 sg13g2_dlygate4sd3_1
Xhold1072 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[6\]
+ VPWR VGND net2899 sg13g2_dlygate4sd3_1
XFILLER_26_84 VPWR VGND sg13g2_fill_1
XFILLER_26_471 VPWR VGND sg13g2_fill_2
XFILLER_53_290 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_117_clk_regs clknet_5_19__leaf_clk_regs clknet_leaf_117_clk_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_42_61 VPWR VGND sg13g2_fill_2
XFILLER_6_821 VPWR VGND sg13g2_fill_1
XFILLER_6_843 VPWR VGND sg13g2_decap_8
XFILLER_5_320 VPWR VGND sg13g2_fill_2
X_08538__142 VPWR VGND net142 sg13g2_tiehi
X_08722__1266 VPWR VGND net1686 sg13g2_tiehi
XFILLER_97_1024 VPWR VGND sg13g2_decap_4
XFILLER_3_1028 VPWR VGND sg13g2_fill_1
X_05620_ net1119 i_exotiny._1924_\[5\] _02286_ VPWR VGND sg13g2_nor2b_1
X_05551_ _02235_ net2735 net1071 VPWR VGND sg13g2_nand2_1
X_08944__1038 VPWR VGND net1458 sg13g2_tiehi
X_08270_ net408 VGND VPWR _00351_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[29\].i_reg.reg_r\[4\]
+ clknet_leaf_101_clk_regs sg13g2_dfrbpq_1
X_05482_ _02182_ net1284 net3584 VPWR VGND sg13g2_nand2_1
XFILLER_32_452 VPWR VGND sg13g2_fill_1
X_07221_ _02971_ VPWR _00946_ VGND _01417_ net1086 sg13g2_o21ai_1
XFILLER_73_0 VPWR VGND sg13g2_fill_2
X_07152_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[13\]
+ net2828 net1009 _00900_ VPWR VGND sg13g2_mux2_1
X_06103_ net2276 _02521_ net957 _00278_ VPWR VGND sg13g2_mux2_1
XFILLER_105_207 VPWR VGND sg13g2_decap_8
X_07083_ net2644 net3404 net915 _00838_ VPWR VGND sg13g2_mux2_1
XFILLER_99_430 VPWR VGND sg13g2_decap_8
X_06034_ net2562 net2521 net962 _00219_ VPWR VGND sg13g2_mux2_1
XFILLER_102_958 VPWR VGND sg13g2_decap_8
XFILLER_101_457 VPWR VGND sg13g2_decap_8
X_07985_ net126 VGND VPWR net2126 i_exotiny._0369_\[9\] clknet_leaf_14_clk_regs sg13g2_dfrbpq_1
X_06936_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[25\].i_reg.reg_r\[16\]
+ net3032 net926 _00715_ VPWR VGND sg13g2_mux2_1
X_06867_ net3620 net1095 _02877_ VPWR VGND sg13g2_nor2_1
XFILLER_103_67 VPWR VGND sg13g2_fill_1
X_05818_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[14\]
+ net2598 net1057 _00090_ VPWR VGND sg13g2_mux2_1
X_08606_ net1790 VGND VPWR net3631 i_exotiny._1614_\[2\] clknet_leaf_23_clk_regs sg13g2_dfrbpq_2
XFILLER_43_706 VPWR VGND sg13g2_decap_8
XFILLER_103_78 VPWR VGND sg13g2_fill_2
X_06798_ VGND VPWR _02816_ _02818_ _02819_ net1130 sg13g2_a21oi_1
X_05749_ net3606 _01584_ _02384_ VPWR VGND sg13g2_nor2_1
X_08537_ net143 VGND VPWR net2151 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[25\]
+ clknet_leaf_183_clk_regs sg13g2_dfrbpq_1
XFILLER_23_441 VPWR VGND sg13g2_fill_2
X_08468_ net212 VGND VPWR net3069 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[20\]
+ clknet_leaf_64_clk_regs sg13g2_dfrbpq_1
XFILLER_23_485 VPWR VGND sg13g2_fill_1
X_07419_ net1082 net2077 _03066_ _01049_ VPWR VGND sg13g2_a21o_1
X_08399_ net683 VGND VPWR net3562 i_exotiny.i_wb_spi.cnt_presc_r\[5\] clknet_leaf_31_clk_regs
+ sg13g2_dfrbpq_1
X_08800__1188 VPWR VGND net1608 sg13g2_tiehi
XFILLER_3_802 VPWR VGND sg13g2_decap_8
XFILLER_88_24 VPWR VGND sg13g2_fill_1
X_08175__502 VPWR VGND net502 sg13g2_tiehi
XFILLER_105_741 VPWR VGND sg13g2_decap_8
Xhold180 _00035_ VPWR VGND net2007 sg13g2_dlygate4sd3_1
XFILLER_3_879 VPWR VGND sg13g2_decap_8
Xhold191 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[23\]
+ VPWR VGND net2018 sg13g2_dlygate4sd3_1
X_09205__776 VPWR VGND net776 sg13g2_tiehi
XFILLER_65_308 VPWR VGND sg13g2_fill_1
XFILLER_59_861 VPWR VGND sg13g2_fill_2
X_08288__390 VPWR VGND net390 sg13g2_tiehi
XFILLER_33_227 VPWR VGND sg13g2_fill_2
XFILLER_61_547 VPWR VGND sg13g2_fill_2
XFILLER_15_953 VPWR VGND sg13g2_fill_2
XFILLER_26_290 VPWR VGND sg13g2_fill_2
XFILLER_15_986 VPWR VGND sg13g2_fill_2
XFILLER_105_1028 VPWR VGND sg13g2_fill_1
X_09112__870 VPWR VGND net870 sg13g2_tiehi
XFILLER_97_912 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_85_clk_regs clknet_5_30__leaf_clk_regs clknet_leaf_85_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08295__383 VPWR VGND net383 sg13g2_tiehi
XFILLER_45_4 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_14_clk_regs clknet_5_6__leaf_clk_regs clknet_leaf_14_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_96_444 VPWR VGND sg13g2_decap_4
Xhold1808 _00859_ VPWR VGND net3635 sg13g2_dlygate4sd3_1
XFILLER_97_989 VPWR VGND sg13g2_decap_8
X_07770_ net2132 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[22\]
+ net988 _01255_ VPWR VGND sg13g2_mux2_1
Xhold1819 i_exotiny.i_wb_spi.dat_rx_r\[29\] VPWR VGND net3646 sg13g2_dlygate4sd3_1
X_04982_ _01712_ _01713_ _01714_ VPWR VGND sg13g2_nor2_1
X_06721_ VGND VPWR _01403_ net1187 _02754_ _02753_ sg13g2_a21oi_1
X_06652_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_wden.u_bit_field.i_sw_write_data[0]
+ _02691_ _02693_ VPWR VGND sg13g2_nor2_1
X_05603_ net1072 _02272_ _02273_ VPWR VGND sg13g2_nor2_1
X_06583_ i_exotiny._0314_\[7\] net1164 _02645_ VPWR VGND sg13g2_nor2_1
X_08322_ net356 VGND VPWR _00403_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[24\]
+ clknet_leaf_83_clk_regs sg13g2_dfrbpq_1
X_05534_ VGND VPWR i_exotiny.i_wb_qspi_mem.crm_r _01520_ _02221_ _01512_ sg13g2_a21oi_1
X_08253_ net424 VGND VPWR _00334_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[24\].i_reg.reg_r\[20\]
+ clknet_leaf_49_clk_regs sg13g2_dfrbpq_1
XFILLER_60_580 VPWR VGND sg13g2_decap_4
XFILLER_32_271 VPWR VGND sg13g2_fill_2
X_07204_ _02964_ net1933 net1088 VPWR VGND sg13g2_nand2_1
X_05465_ _02171_ _02149_ i_exotiny._1617_\[3\] _02148_ i_exotiny._1612_\[3\] VPWR
+ VGND sg13g2_a22oi_1
X_05396_ net1112 _02112_ i_exotiny._2043_\[2\] VPWR VGND sg13g2_nor2_1
X_08184_ net493 VGND VPWR net2074 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[4\].i_reg.reg_r\[15\]
+ clknet_leaf_109_clk_regs sg13g2_dfrbpq_1
X_07981__122 VPWR VGND net122 sg13g2_tiehi
X_07135_ net1286 net1834 _00885_ VPWR VGND sg13g2_and2_1
XFILLER_106_538 VPWR VGND sg13g2_decap_8
X_07066_ net2866 net878 _02934_ _02938_ VPWR VGND sg13g2_mux2_1
X_08159__519 VPWR VGND net519 sg13g2_tiehi
X_06017_ _00018_ net1103 _02503_ VPWR VGND sg13g2_nor2_1
XFILLER_0_805 VPWR VGND sg13g2_decap_8
XFILLER_102_766 VPWR VGND sg13g2_fill_1
XFILLER_101_254 VPWR VGND sg13g2_decap_8
X_07968_ net1177 VGND VPWR net3793 i_exotiny.i_wdg_top.o_wb_dat\[9\] clknet_leaf_35_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_68_691 VPWR VGND sg13g2_fill_1
X_06919_ _02916_ net1138 net1165 _02917_ VPWR VGND sg13g2_a21o_2
X_07899_ net45 VGND VPWR _00001_ i_exotiny._1312_ clknet_leaf_13_clk_regs sg13g2_dfrbpq_1
X_08528__152 VPWR VGND net152 sg13g2_tiehi
XFILLER_70_333 VPWR VGND sg13g2_fill_1
XFILLER_51_591 VPWR VGND sg13g2_fill_2
XFILLER_8_916 VPWR VGND sg13g2_decap_8
XFILLER_12_967 VPWR VGND sg13g2_decap_8
XFILLER_23_293 VPWR VGND sg13g2_fill_1
X_08396__536 VPWR VGND net536 sg13g2_tiehi
X_08535__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_105_571 VPWR VGND sg13g2_decap_8
XFILLER_79_945 VPWR VGND sg13g2_fill_2
XFILLER_94_948 VPWR VGND sg13g2_decap_8
XFILLER_17_8 VPWR VGND sg13g2_decap_4
XFILLER_47_875 VPWR VGND sg13g2_fill_1
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_34_525 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_132_clk_regs clknet_5_20__leaf_clk_regs clknet_leaf_132_clk_regs VPWR
+ VGND sg13g2_buf_8
X_08542__138 VPWR VGND net138 sg13g2_tiehi
XFILLER_9_32 VPWR VGND sg13g2_fill_2
XFILLER_9_76 VPWR VGND sg13g2_fill_1
X_05250_ _01831_ VPWR _01976_ VGND _01974_ _01975_ sg13g2_o21ai_1
X_05181_ _01900_ _01904_ _01906_ _01909_ VPWR VGND sg13g2_nor3_1
Xhold916 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[15\]
+ VPWR VGND net2743 sg13g2_dlygate4sd3_1
Xhold905 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[27\]
+ VPWR VGND net2732 sg13g2_dlygate4sd3_1
Xhold927 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[24\]
+ VPWR VGND net2754 sg13g2_dlygate4sd3_1
XFILLER_7_982 VPWR VGND sg13g2_decap_8
Xhold949 _00421_ VPWR VGND net2776 sg13g2_dlygate4sd3_1
Xhold938 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[28\].i_reg.reg_r\[8\]
+ VPWR VGND net2765 sg13g2_dlygate4sd3_1
X_08940_ net1462 VGND VPWR net2585 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[6\]
+ clknet_leaf_74_clk_regs sg13g2_dfrbpq_1
X_08894__1088 VPWR VGND net1508 sg13g2_tiehi
X_08871_ net1531 VGND VPWR net3590 i_exotiny.i_wb_spi.dat_rx_r\[1\] clknet_leaf_28_clk_regs
+ sg13g2_dfrbpq_1
XFILLER_9_1023 VPWR VGND sg13g2_decap_4
X_08582__1398 VPWR VGND net1818 sg13g2_tiehi
XFILLER_36_0 VPWR VGND sg13g2_decap_8
Xhold1605 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[16\]
+ VPWR VGND net3432 sg13g2_dlygate4sd3_1
Xhold1616 i_exotiny._0369_\[10\] VPWR VGND net3443 sg13g2_dlygate4sd3_1
X_07822_ _02477_ _02525_ _03222_ VPWR VGND sg13g2_nor2_2
Xhold1627 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[19\]
+ VPWR VGND net3454 sg13g2_dlygate4sd3_1
Xhold1649 i_exotiny._0314_\[8\] VPWR VGND net3476 sg13g2_dlygate4sd3_1
Xhold1638 _00853_ VPWR VGND net3465 sg13g2_dlygate4sd3_1
X_07753_ net2900 net2600 net991 _01238_ VPWR VGND sg13g2_mux2_1
XFILLER_38_875 VPWR VGND sg13g2_fill_2
X_04965_ _01697_ _01362_ _01696_ VPWR VGND sg13g2_nand2b_1
XFILLER_93_970 VPWR VGND sg13g2_decap_8
X_06704_ _02739_ i_exotiny.gpo\[2\] _02725_ VPWR VGND sg13g2_nand2_1
X_07684_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[19\]
+ net2176 net998 _01186_ VPWR VGND sg13g2_mux2_1
X_04896_ i_exotiny._0077_\[2\] i_exotiny._0077_\[3\] net1257 _01628_ VGND VPWR _01617_
+ sg13g2_nor4_2
X_06635_ net2446 net1152 _02680_ VPWR VGND sg13g2_nor2_1
XFILLER_12_208 VPWR VGND sg13g2_fill_2
X_08305_ net373 VGND VPWR _00386_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[27\].i_reg.reg_r\[7\]
+ clknet_leaf_73_clk_regs sg13g2_dfrbpq_1
X_06566_ net3603 net1154 _02634_ VPWR VGND sg13g2_nor2_1
X_06497_ net2561 net2228 net1026 _00578_ VPWR VGND sg13g2_mux2_1
X_09285_ net51 VGND VPWR net2189 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[18\].i_reg.reg_r\[11\]
+ clknet_leaf_168_clk_regs sg13g2_dfrbpq_1
X_05517_ VGND VPWR i_exotiny._0314_\[11\] net1276 _02208_ _02207_ sg13g2_a21oi_1
X_08236_ net441 VGND VPWR net3103 i_exotiny._0028_\[3\] clknet_leaf_60_clk_regs sg13g2_dfrbpq_2
X_05448_ _02156_ _02140_ i_exotiny._1618_\[1\] _02135_ i_exotiny._1614_\[1\] VPWR
+ VGND sg13g2_a22oi_1
X_08681__1307 VPWR VGND net1727 sg13g2_tiehi
X_08167_ net511 VGND VPWR net2801 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[31\]
+ clknet_leaf_119_clk_regs sg13g2_dfrbpq_1
X_07118_ net1288 net1847 _00868_ VPWR VGND sg13g2_and2_1
X_05379_ i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_hw_set[0]
+ net3780 _02076_ _02101_ VPWR VGND sg13g2_nor3_1
XFILLER_106_335 VPWR VGND sg13g2_decap_8
X_08098_ net596 VGND VPWR _00179_ i_exotiny._0013_\[3\] clknet_leaf_125_clk_regs sg13g2_dfrbpq_2
X_07049_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[19\]
+ net3199 net1016 _00810_ VPWR VGND sg13g2_mux2_1
XFILLER_88_720 VPWR VGND sg13g2_fill_1
X_08172__505 VPWR VGND net505 sg13g2_tiehi
XFILLER_102_541 VPWR VGND sg13g2_fill_2
XFILLER_102_574 VPWR VGND sg13g2_fill_2
XFILLER_47_105 VPWR VGND sg13g2_fill_1
X_09202__779 VPWR VGND net779 sg13g2_tiehi
X_09102__880 VPWR VGND net1300 sg13g2_tiehi
Xclkbuf_5_15__f_clk_regs clknet_4_7_0_clk_regs clknet_5_15__leaf_clk_regs VPWR VGND
+ sg13g2_buf_8
XFILLER_55_182 VPWR VGND sg13g2_fill_2
XFILLER_16_536 VPWR VGND sg13g2_fill_2
X_08285__393 VPWR VGND net393 sg13g2_tiehi
X_08657__1320 VPWR VGND net1740 sg13g2_tiehi
XFILLER_4_974 VPWR VGND sg13g2_decap_8
XFILLER_78_263 VPWR VGND sg13g2_fill_2
X_08292__386 VPWR VGND net386 sg13g2_tiehi
Xfanout1230 net3699 net1230 VPWR VGND sg13g2_buf_8
Xfanout1241 net3837 net1241 VPWR VGND sg13g2_buf_2
Xfanout1263 i_exotiny.i_wdg_top.wdgrv_regs_inst.g_wdcsr.g_s1wto.u_bit_field.i_hw_set[0]
+ net1263 VPWR VGND sg13g2_buf_8
Xfanout1274 i_exotiny._1312_ net1274 VPWR VGND sg13g2_buf_8
Xfanout1252 i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.i_r\[3\]
+ net1252 VPWR VGND sg13g2_buf_8
Xfanout1285 net1291 net1285 VPWR VGND sg13g2_buf_8
X_08879__1103 VPWR VGND net1523 sg13g2_tiehi
X_04750_ _01504_ net1279 net3705 VPWR VGND sg13g2_nand2_1
XFILLER_90_940 VPWR VGND sg13g2_decap_8
XFILLER_74_480 VPWR VGND sg13g2_decap_8
XFILLER_62_631 VPWR VGND sg13g2_fill_1
X_06420_ net3730 _02595_ _02600_ VPWR VGND sg13g2_nor2_1
X_08149__529 VPWR VGND net529 sg13g2_tiehi
X_04681_ _01441_ VPWR i_exotiny._1489_\[3\] VGND net1266 _01438_ sg13g2_o21ai_1
X_06351_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[30\].i_reg.reg_r\[10\]
+ net3373 net1030 _00481_ VPWR VGND sg13g2_mux2_1
X_09070_ net1332 VGND VPWR net1879 i_exotiny.i_wdg_top.clk_div_inst.cnt\[10\] clknet_leaf_45_clk_regs
+ sg13g2_dfrbpq_1
X_06282_ net2963 net2775 net944 _00425_ VPWR VGND sg13g2_mux2_1
X_05302_ _02028_ _01655_ i_exotiny._0026_\[0\] _01651_ i_exotiny._0039_\[0\] VPWR
+ VGND sg13g2_a22oi_1
X_08021_ net673 VGND VPWR _00102_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[22\]
+ clknet_leaf_61_clk_regs sg13g2_dfrbpq_1
X_05233_ _01961_ _01630_ i_exotiny._0041_\[1\] _01619_ i_exotiny._0034_\[1\] VPWR
+ VGND sg13g2_a22oi_1
Xhold702 _00049_ VPWR VGND net2529 sg13g2_dlygate4sd3_1
Xhold746 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[21\]
+ VPWR VGND net2573 sg13g2_dlygate4sd3_1
Xhold713 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[11\]
+ VPWR VGND net2540 sg13g2_dlygate4sd3_1
Xhold724 _00532_ VPWR VGND net2551 sg13g2_dlygate4sd3_1
XFILLER_7_790 VPWR VGND sg13g2_decap_4
Xhold735 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[21\].i_reg.reg_r\[6\]
+ VPWR VGND net2562 sg13g2_dlygate4sd3_1
X_05164_ _01880_ _01883_ _01879_ _01894_ VPWR VGND _01893_ sg13g2_nand4_1
XFILLER_104_839 VPWR VGND sg13g2_decap_8
Xhold757 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[10\]
+ VPWR VGND net2584 sg13g2_dlygate4sd3_1
Xhold779 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[9\].i_reg.reg_r\[15\]
+ VPWR VGND net2606 sg13g2_dlygate4sd3_1
X_08518__162 VPWR VGND net162 sg13g2_tiehi
X_05095_ VPWR VGND _01814_ net1110 _01752_ i_exotiny.i_fazyrv_top.i_fazyrv_core.genblk2.i_fazyrv_decode.imm_o\[3\]
+ _01826_ net1108 sg13g2_a221oi_1
Xhold768 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[13\]
+ VPWR VGND net2595 sg13g2_dlygate4sd3_1
X_08923_ net1479 VGND VPWR net2714 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[21\]
+ clknet_leaf_113_clk_regs sg13g2_dfrbpq_1
XFILLER_39_18 VPWR VGND sg13g2_fill_1
Xhold1402 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[13\].i_reg.reg_r\[26\]
+ VPWR VGND net3229 sg13g2_dlygate4sd3_1
X_08854_ net1552 VGND VPWR _00912_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[21\]
+ clknet_leaf_186_clk_regs sg13g2_dfrbpq_1
Xhold1424 _01343_ VPWR VGND net3251 sg13g2_dlygate4sd3_1
Xhold1413 _00616_ VPWR VGND net3240 sg13g2_dlygate4sd3_1
Xhold1468 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[10\]
+ VPWR VGND net3295 sg13g2_dlygate4sd3_1
Xhold1457 _00160_ VPWR VGND net3284 sg13g2_dlygate4sd3_1
Xhold1435 _00480_ VPWR VGND net3262 sg13g2_dlygate4sd3_1
X_07805_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[1\].i_reg.reg_r\[19\]
+ net2345 net891 _01284_ VPWR VGND sg13g2_mux2_1
X_08785_ net1623 VGND VPWR net2968 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[16\]
+ clknet_leaf_167_clk_regs sg13g2_dfrbpq_1
Xhold1446 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[25\]
+ VPWR VGND net3273 sg13g2_dlygate4sd3_1
X_05997_ net2337 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[27\]
+ net1051 _00199_ VPWR VGND sg13g2_mux2_1
Xhold1479 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[28\]
+ VPWR VGND net3306 sg13g2_dlygate4sd3_1
X_07736_ _03203_ net2517 net996 _01229_ VPWR VGND sg13g2_mux2_1
X_04948_ net1242 _01533_ _01604_ _01680_ VPWR VGND sg13g2_nor3_1
X_08735__1253 VPWR VGND net1673 sg13g2_tiehi
X_08525__155 VPWR VGND net155 sg13g2_tiehi
XFILLER_25_355 VPWR VGND sg13g2_fill_1
X_07667_ net2511 net2899 net1001 _01169_ VPWR VGND sg13g2_mux2_1
X_04879_ _01611_ _01460_ _01602_ _01421_ net1254 VPWR VGND sg13g2_a22oi_1
X_07598_ _03170_ i_exotiny.i_wdg_top.clk_div_inst.cnt\[9\] net1877 _03166_ VPWR VGND
+ sg13g2_and3_2
XFILLER_52_185 VPWR VGND sg13g2_fill_1
XFILLER_52_163 VPWR VGND sg13g2_fill_1
X_06618_ net1199 _02667_ _02668_ _00646_ VPWR VGND sg13g2_nor3_1
X_06549_ net1210 net3757 _02626_ _00619_ VPWR VGND sg13g2_a21o_1
X_09268_ net91 VGND VPWR net2122 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[26\]
+ clknet_leaf_127_clk_regs sg13g2_dfrbpq_1
X_08219_ net458 VGND VPWR net2262 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[3\].i_reg.reg_r\[18\]
+ clknet_leaf_151_clk_regs sg13g2_dfrbpq_1
X_09199_ net782 VGND VPWR _01254_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[22\].i_reg.reg_r\[21\]
+ clknet_leaf_78_clk_regs sg13g2_dfrbpq_1
XFILLER_106_132 VPWR VGND sg13g2_decap_8
X_08957__1025 VPWR VGND net1445 sg13g2_tiehi
X_08532__148 VPWR VGND net148 sg13g2_tiehi
XFILLER_1_922 VPWR VGND sg13g2_decap_8
XFILLER_0_454 VPWR VGND sg13g2_fill_1
XFILLER_102_371 VPWR VGND sg13g2_decap_8
Xhold40 i_exotiny.i_wb_spi.state_r\[16\] VPWR VGND net1867 sg13g2_dlygate4sd3_1
XFILLER_0_465 VPWR VGND sg13g2_fill_2
XFILLER_1_999 VPWR VGND sg13g2_decap_8
Xhold51 _03169_ VPWR VGND net1878 sg13g2_dlygate4sd3_1
Xhold62 _00076_ VPWR VGND net1889 sg13g2_dlygate4sd3_1
Xhold73 _00054_ VPWR VGND net1900 sg13g2_dlygate4sd3_1
XFILLER_91_715 VPWR VGND sg13g2_fill_2
Xhold95 i_exotiny._1924_\[12\] VPWR VGND net1922 sg13g2_dlygate4sd3_1
Xhold84 i_exotiny._1160_\[27\] VPWR VGND net1911 sg13g2_dlygate4sd3_1
Xhold1980 i_exotiny._0542_ VPWR VGND net3807 sg13g2_dlygate4sd3_1
XFILLER_16_311 VPWR VGND sg13g2_fill_2
Xhold1991 i_exotiny._0077_\[3\] VPWR VGND net3818 sg13g2_dlygate4sd3_1
XFILLER_91_1008 VPWR VGND sg13g2_decap_8
X_08867__1118 VPWR VGND net1538 sg13g2_tiehi
XFILLER_16_366 VPWR VGND sg13g2_fill_1
XFILLER_44_653 VPWR VGND sg13g2_fill_2
XFILLER_31_314 VPWR VGND sg13g2_fill_1
X_08606__1370 VPWR VGND net1790 sg13g2_tiehi
XFILLER_4_771 VPWR VGND sg13g2_decap_8
X_08813__1175 VPWR VGND net1595 sg13g2_tiehi
XFILLER_98_369 VPWR VGND sg13g2_decap_8
X_05920_ net2164 net2444 net972 _00137_ VPWR VGND sg13g2_mux2_1
XFILLER_6_1004 VPWR VGND sg13g2_decap_8
XFILLER_94_542 VPWR VGND sg13g2_fill_1
Xfanout1060 net1061 net1060 VPWR VGND sg13g2_buf_1
X_05851_ _02439_ VPWR _02440_ VGND _02055_ _02069_ sg13g2_o21ai_1
Xfanout1082 net1084 net1082 VPWR VGND sg13g2_buf_8
Xfanout1071 _02181_ net1071 VPWR VGND sg13g2_buf_8
XFILLER_94_597 VPWR VGND sg13g2_fill_1
X_04802_ VGND VPWR _01549_ _01548_ i_exotiny._3871_ sg13g2_or2_1
Xfanout1093 _02960_ net1093 VPWR VGND sg13g2_buf_8
X_08570_ net64 VGND VPWR net3244 i_exotiny._0314_\[15\] clknet_leaf_180_clk_regs sg13g2_dfrbpq_1
X_05782_ net3715 VPWR _00073_ VGND net1143 _02404_ sg13g2_o21ai_1
X_07521_ net901 net3570 _03118_ _01099_ VPWR VGND sg13g2_a21o_1
Xclkbuf_4_12_0_clk_regs clknet_0_clk_regs clknet_4_12_0_clk_regs VPWR VGND sg13g2_buf_8
X_04733_ i_exotiny._0315_\[28\] i_exotiny._0314_\[28\] net1271 _01489_ VPWR VGND sg13g2_mux2_1
XFILLER_62_472 VPWR VGND sg13g2_fill_2
X_04664_ _01425_ _01420_ _01423_ VPWR VGND sg13g2_nand2_2
X_07452_ VGND VPWR net3535 net1080 _03091_ _03077_ sg13g2_a21oi_1
XFILLER_23_859 VPWR VGND sg13g2_fill_1
X_06403_ _02587_ _02586_ _01512_ _01520_ _01485_ VPWR VGND sg13g2_a22oi_1
X_07383_ _03038_ _03025_ _03037_ net1210 i_exotiny._1160_\[9\] VPWR VGND sg13g2_a22oi_1
X_06334_ net3260 net887 _02558_ _02560_ VPWR VGND sg13g2_mux2_1
X_09122_ net860 VGND VPWR _01177_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[26\].i_reg.reg_r\[10\]
+ clknet_leaf_157_clk_regs sg13g2_dfrbpq_1
X_09053_ net1349 VGND VPWR _01108_ i_exotiny.i_rstctl.cnt\[3\] clknet_leaf_39_clk_regs
+ sg13g2_dfrbpq_1
X_06265_ _02551_ net2640 net1039 _00410_ VPWR VGND sg13g2_mux2_1
X_08004_ net691 VGND VPWR net2322 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[15\].i_reg.reg_r\[5\]
+ clknet_leaf_66_clk_regs sg13g2_dfrbpq_1
X_06196_ net2629 net2146 net948 _00351_ VPWR VGND sg13g2_mux2_1
X_05216_ VGND VPWR _01750_ _01943_ _01944_ net1108 sg13g2_a21oi_1
Xhold510 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[10\].i_reg.reg_r\[23\]
+ VPWR VGND net2337 sg13g2_dlygate4sd3_1
Xhold543 _00368_ VPWR VGND net2370 sg13g2_dlygate4sd3_1
Xhold521 _01318_ VPWR VGND net2348 sg13g2_dlygate4sd3_1
Xhold532 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[12\].i_reg.reg_r\[7\]
+ VPWR VGND net2359 sg13g2_dlygate4sd3_1
Xhold554 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[17\]
+ VPWR VGND net2381 sg13g2_dlygate4sd3_1
X_05147_ _01877_ _01646_ i_exotiny._0017_\[2\] _01632_ i_exotiny._0022_\[2\] VPWR
+ VGND sg13g2_a22oi_1
Xhold587 _00268_ VPWR VGND net2414 sg13g2_dlygate4sd3_1
Xhold576 _00415_ VPWR VGND net2403 sg13g2_dlygate4sd3_1
Xhold565 _00238_ VPWR VGND net2392 sg13g2_dlygate4sd3_1
XFILLER_106_45 VPWR VGND sg13g2_fill_2
XFILLER_103_157 VPWR VGND sg13g2_decap_8
XFILLER_89_358 VPWR VGND sg13g2_fill_2
Xhold598 _00440_ VPWR VGND net2425 sg13g2_dlygate4sd3_1
X_05078_ _01808_ _01809_ _01807_ _01810_ VPWR VGND sg13g2_nand3_1
XFILLER_98_881 VPWR VGND sg13g2_decap_8
XFILLER_97_380 VPWR VGND sg13g2_decap_8
X_08906_ net1496 VGND VPWR net3315 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[6\].i_reg.reg_r\[4\]
+ clknet_leaf_65_clk_regs sg13g2_dfrbpq_1
Xhold1232 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[8\].i_reg.reg_r\[26\]
+ VPWR VGND net3059 sg13g2_dlygate4sd3_1
Xhold1243 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[20\].i_reg.reg_r\[23\]
+ VPWR VGND net3070 sg13g2_dlygate4sd3_1
X_08837_ net1569 VGND VPWR _00895_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[31\].i_reg.reg_r\[4\]
+ clknet_leaf_184_clk_regs sg13g2_dfrbpq_1
Xhold1210 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[5\].i_reg.reg_r\[5\]
+ VPWR VGND net3037 sg13g2_dlygate4sd3_1
Xhold1221 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[19\].i_reg.reg_r\[10\]
+ VPWR VGND net3048 sg13g2_dlygate4sd3_1
XFILLER_100_875 VPWR VGND sg13g2_decap_8
Xhold1265 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[16\].i_reg.reg_r\[8\]
+ VPWR VGND net3092 sg13g2_dlygate4sd3_1
Xhold1254 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[17\].i_reg.reg_r\[7\]
+ VPWR VGND net3081 sg13g2_dlygate4sd3_1
Xhold1276 _00317_ VPWR VGND net3103 sg13g2_dlygate4sd3_1
X_08768_ net1640 VGND VPWR _00826_ i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[14\].i_reg.reg_r\[31\]
+ clknet_leaf_81_clk_regs sg13g2_dfrbpq_1
Xhold1287 _01092_ VPWR VGND net3114 sg13g2_dlygate4sd3_1
Xhold1298 _01302_ VPWR VGND net3125 sg13g2_dlygate4sd3_1
X_08699_ net1709 VGND VPWR net2161 i_exotiny.i_fazyrv_top.genblk2.i_fazyrv_rf_lut.genblk1\[2\].i_reg.reg_r\[26\]
+ clknet_leaf_105_clk_regs sg13g2_dfrbpq_1
X_07719_ net3090 net2916 net993 _01215_ VPWR VGND sg13g2_mux2_1
X_08282__396 VPWR VGND net396 sg13g2_tiehi
XFILLER_12_1009 VPWR VGND sg13g2_decap_8
XFILLER_5_513 VPWR VGND sg13g2_fill_2
XFILLER_103_0 VPWR VGND sg13g2_fill_2
Xoutput41 net41 uo_out[7] VPWR VGND sg13g2_buf_1
Xoutput30 net30 uio_out[4] VPWR VGND sg13g2_buf_1
XFILLER_95_328 VPWR VGND sg13g2_decap_8
XFILLER_49_701 VPWR VGND sg13g2_fill_2
XFILLER_1_796 VPWR VGND sg13g2_decap_8
XFILLER_49_789 VPWR VGND sg13g2_fill_2
XFILLER_17_631 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_39_clk_regs clknet_5_10__leaf_clk_regs clknet_leaf_39_clk_regs VPWR VGND
+ sg13g2_buf_8
X_08508__172 VPWR VGND net172 sg13g2_tiehi
XFILLER_32_612 VPWR VGND sg13g2_fill_2
XFILLER_16_196 VPWR VGND sg13g2_fill_2
X_06050_ net2699 net3025 net961 _00235_ VPWR VGND sg13g2_mux2_1
X_05001_ net1174 _01705_ _01724_ _01733_ VPWR VGND sg13g2_nor3_1
XFILLER_59_509 VPWR VGND sg13g2_decap_4
X_08515__165 VPWR VGND net165 sg13g2_tiehi
X_06952_ net3043 net877 _02916_ _02920_ VPWR VGND sg13g2_mux2_1
.ends

