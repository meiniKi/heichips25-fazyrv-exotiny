`default_nettype none

module fazyrv_small_logo ();
endmodule
